��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su˸Y��'��d�Ay~�`�i���o3 1&����1\T�����	��!mF��
��\�ݘ�#X4|'�~a	N�1�""rϗ��?���ݝ��^��lt����d�k>O@�0�#/���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�Oo�Ne�<��!G�u�uO]�nG����W��1L���a�KzܸƠC[#f�0�����-V_� 8T^(�|��Z0��+����[VT`�c��A�p�����	�S��60�W���)/��L��A�g87V�c�5�_Җ��sd�����PA��C%#!^��M[��[C�r��O�k�#H�w�c���T��7rC��i ��)�sI?�V�K7ۉ0���F4rg���W��:����J����Em��]������ \do<<(���1�'��*��{�"�%4P�D��V"R��G�xVxV����\��T:r/����q�B3�z��2z��un/D��QG%�=oTK�;�I%�ǿ���α��|��mی���o������?��H��t�x��M���ug"A��w� ��fS��������`���?��X���N�����^T(�u��p������l�YA?����L��bI���7lc�f�6FnEq��Fl��� ��g�Y�)RyX蚞�u����^�vTC��n���S���]���TWq�x�B��˽{��`��*����h*CN@�-�C>�_i���8_DyS�b�ʥ�^vo�0w�����a�?�1n� ��Ǭ� AR�ϓ\6��bu�_"[�P8p���	��1� �өVt� .m3�p���Qr�%���Z�^��'VHDb
v4�;/��u�_��e�T�ÙRj��]���u]/GR�r�ۣ|w{拈�?��x�N-�,����=����B�H
�b^"�׉��i���+$}\T~YַD�K�1B��q����u�(Rc{3=����ng�8Z���5� ṘB��h��T<�;92��W���}������F�b�I�:y><��#�c���Vn4�{Ʀ1��Qx�b*�G	� ��5_�����քl��l4���e�Iݞ>�#6A���ؼ=�gi��6	���D�8�/Y�ėגZu'���^��YD 0�^��q�<�l�Ϻ��+z���L#�ʦ�LA���d���t�.�PT4"�̣�H!J�5G���zR��h�x���2�E:�X������Ѻth7�]\r��cqc�\����.o��g�fC�D���	,�sg�P&�˸������p���s/ǱB6����zNz�RGjӻt5�E�8(�Յ�+8����!��[�ݦ�m���HI�_��.~�\���X�`��~!�j�M�u�O�!��:�%g|0�c�P��?p�O�>T��(��1�K%�Bsvs�8��d���Ë��43�P���9�0�?�����6��o�E�|�,�ER Af#/y�lY�B���GK���ڒ�GBR@$<3�F4�8E�6]��͢Y��"ܾ�T�ݧ��bP"ְb�5f�:|����)*�>�&E"�-����J�)zVi�?��{�p�3���F�&I���ح���h� <A����r(?%2�vZK�!�ԑ���� �z��f+�gvaGֳ����7��	)����;L�nx���7�c�e�DE`0����Y�Wkjv䬒�4��l�~�]3��(��>*��G��B����b%�𝬟n�,*`��M����W�������_
��s>��~ ��swq�^ޑ�L�]���s��Bl�x�;F�g��yۿ�Y����ڔ�"�F�+��o�_=��:.Ȫ7	�>�z����Ò���r�jcX��XK�%uső������o�+�����?����H}-��sL�idX/�[o*�AjK��UvFؚI�nj8䠮���/y>�����O�&	�H^�p)�
\
�j��
�b�i�<[��3�ݸ�4My��f�K���~Y���X��r�]?�C�N�ä���Κ��:2��O�JF{���W[r�(�����_�"��� �=�7�eX�X�&A��ߏW,�/���<ϊz7f���N��1����|{&��V6>A�C�vAYq([����Il�cZjٶ�I�x�tBi�ISi����eM.��%p-�N��kAz�/�1*�߅����r�|��5��v���&=�O�.�E: gX�TK4����Q�d?|�D_ � �� G~�{ڝO��#0�K�,��Zd\oB�&�`��O��Qf�:�� o�+E�����H{ŕ �DC>��P������Fg�q����� ���Q�3(|S)����SZ36q�zc}^V8�"V�'�r~�q�KB}A�����)9�y�yXVR� ��ָ��m���N����@��S���q:J�(������8F~��E���G������c,8��:E/����WPh���i��7�Wi��������q���e��p��X)��p	��O4P��n�0x��` Rҿ�
>%�'��&�ڝmNqb��;]�NPz�1�	Sp��,}V�BqJЗa�b@�;���k ���dOo�n�]� �i��W��X7�)%Ok�S�E���E���<h;��ץ�|�O��h���ށ?���#�� C�{���lբ�!ӼN��VW���-l�U3 T�95�Fj�&Ht+D����O�*D!C�n�'t�5պ���=p����������K ��s��n�g{#ofu� �l�v�=I������F/*�g�*x�+��m�0]��5�m���	��j2i�cx_l|;�S��Q�4*a0��]VDi�#�;��ya)q�Ix"��5���[lnx0���t S�`Qv!;^]��G�uC	��~f��<����#��v�l|Q��a�3^Ä��z�d`�X��$�V	�d,ڦ���_J�&|N�<��Nu�C�fi��"g��G��.Z��
kYZ 3,M�����/>�ϸ�)t��U*L|�G�!�ǜN^�"uK.Q��Sw��JGK�PmD�4�DvU^lMZ� �-��4��������ϋJb�K__V����J�_@<���ج��ފOAm7��LBnv�o��JL�Z�?G�K��Jg�Jx����W��]F�����f�G0�#��tx�2��ec��}d.ܖ�ߙ��nɨR �ˑ�Β4���0B�a��_�xW�_j/v�����'	ΞҁN��G�GL2@�L�R;J� r�94�of���3\/`o@:�+M�V��)�a���s$ft�}�O�ў�"*]@��C��`%�ݦOՃ<��A�ͱ0o��/�(�~7�0k���GN��R����!H���Ê��9��C�&v�b�l��c])gY ����O�Voµ���D���%K���u�C0�n�9�c�"�!1��n��s�S�bhopIm���Xа�A
��'zz5���"`c�Çv�7�b��,�^Y���#s@��j�p������I�s��D�&	�P��*�8iP�[�r���y���o�
.�V$T���ף�  C*xJD5�]�/�-����z������lX�c�_T�ŋjVbZ.�NI�,TߵM�[քVv�Ч(
,����p�m`�B7=Y�?Z@�-��g����3
�@x�xt��H�*�5�{ԡ�硵l��{$f��*���nn&��J�Yw(�q;q��BXKG�����a|e,���A��B?�
H�76��t?rzjYm6q�+�3�2��7v|ާ���l�6�`4U]5P��˜�d���9��0av	:�ū9]WfXK`�����xʎI[�(�7�І�$��o2FKҧ"��S<�~|y�a��;�pR�F|�1�ེvY��e*4�{�9���!Uj@K���,��?���U�i��9�X�ѽ�I�y�j�B��[�H��o*�UP��\7���b��2N��I�����Q�9|�U�B��a=��=?�#��K*jWZ�'�+�Մ�3�m<7z����#6������a�D�����tz?it��Ύ�2$
�.<M^BC &�;;w��$5�O����P���sُ'�����:&�j}t��[�_�<�]�AU�S��;22���23~����z��i�ͅw��@�Տ���	�0N���ش9 =`45Kv��I�R����Ol��%�Gإ��(�+��q�%` T�'���+ ��߅�����(�}���2X\=�f�Y�����ǩޏ��GnM�Yof���@I�p+{��LY�v΂r�EP{p�kP�s}���D~�������I5X�b�����(Y����6+o������7�!I���a��p�S��g�e��5aȂ"�iâ�hc<(!��mW�M�r�㠊5��058�i������E��;/1MA������Z�Z�K�K������!���d�/ۺ��|8Wx�d �V�B�L�N(��t�˴3������eu�9�(��������3���6��A�n��1��P��w����V�SM���C+�Z���c4oP\�r���c}]��sx��j4ԁ|IXl���_�6��ޭr8�٨�1dq=KՎ�}X��b��a,�����mE��Z�1�4���ؔg�L�a7�Q��KH<��Sc1����&Hǎ�����/E���I���Q'�S=~�~�����[� �ҽC_�~<��"���%�I������\��	��uڸ���np�Ta��X�M��ȳ��^G�͊Z���Z��l���n*�@��&b"	��)#�}~����hˌr�ԙ�f4E�+|��vR���Z��0E�%C������!�y�^��<Oe��޿}�$�"�/~$4{�w���+CF�R�3/65ޱM�U��%D4�(B��œU#�Q��:���*��ߜV��U�r�PS�'.�}���	'v�.�n�p�#�����E=�韰1M3Sޅ�:h�Wa��^�L��sI�,O�$�ҞE�a����1v�'E0��R��W��ou ��;����+��U=PԽo��u�|��螌��V����'Zo���T���t��67��\�0��O\a���O��8��q�|v2���/}�������OEQN�ؒ�v�4e�=&�^�6.��tn.z�� *��n����ӒT����&` ��<qC��*t$�~0d�Z�Ze��L���B��3B�P��Q��3L��AW���<�PƄ`hd���1�8�J�-�	������)5zO���沥��m1��~T�]�y1�B�t�N��ի��.�R3��D��E�<T�0�2 �/�/LK�����)�} ���/�*[6�����s%�[������� �RF���+0� ļHl,����
��#��%�lx\c��k� �ah��
A�m�p6�I֒)/0��O�D�,*�-�hq�(w!��.^�\_��.F����F��s�nV���i/���g�>(C���妆�.G����3i�f�ɟ��~�g-��cQ ��$_x���ܴ@�d��`l:���4?vW۫N^"#��,�hx��N�f�˸��l�!���+�j�����O�pݚ��ihA���?�LxUt?pZ�x�\�.���N�i6t����cʘ��޷�[��<BA�B�}�us�1�n�vݸ2d	���j=s�ݜ!��QV�0��͗
ϒ�v�M�Rތ��r�w�|�������ES���.�D�ei>)I��P�څ��G��A���ÑHw!.������%��^���;��#��t8��nkV*�OZ�&K:�l&�1WV���,���`t�sӡg3[�A��m����6��:w�X�f�Z�:$��Bȭf��z�x<�Z�<�d��w!��O�" �7��=�A�}Ml3��V��I<V�h��ڨY,����7��\X	�w�4������a��mϔB媲��p3�pyF���R7�ψvR����S2@�����T�A>�&ѣ��m���Q��a;�v�E����Uܙ��\� _#��:&ȋp1*��AT�$ϳ��H��o��(~��|aq��g��X���3BJ�����ڠ�}�F9^�jC��$ejH����L��(�c�*b�#�������|�n|t�sIe���S�&e�5�Ex*�cm�9�e�W\8���I�u7�X�����g	v����%�RgͰɉ�K����$�W���ՁQ��Մ(|3���9��H��nަ��)ݕ�EsTW����g� �3N��cm뿃�(o��@kV�%�;����� �޳�9�����D��ͮ����̔o�e��H�[@[*�nw}^c�_��K��	��������z����׻��v��	����^��@4`�tȤq���vB�lt2���=���GTo�%�|��4[6�� u���Qv�����'����G�:7m'�ޢ�h:;)�<\20�뀲� П��ꊵ����og��TIL�}��:�4H<LB�=�6��9��C�h�0�H�줹0��w�m��W< ���藏ME'��S�������x�v��i$����x/4���^֨�R��h0�J��>"[�`򻧼��E����Ҍں}p!{,8ZC���P�Z��!���f��S������wX=�s���ej�U��'o9�Fs���d���{8`&��oZy_%#�7��i����`���������W����4My��m�0��CB�[�w&�u#����!��	�UR�q�p��]�q�!.QdB�C_�e��H�Y�eY���g}�/\t!����Ę����5���dzp 5f�"���͓��}[	��.������׃S����r�4�.E`d ��*��it0�cn:���T�e_z�#�7�9�%�8P<�ܰq�-��O)4�l_�R �|��������{���s���u$�(��}%VP�� �����7��nqh����3*l%}E��������a�M(�pv�_X����!jGM�5�GP`y�U�����������Ǉ7��덆��RA��7Uiĳ$^ĸޘ\��5#�=UnoG�2?�aH���Aׄ
���'a:�"�;���kV�9��ҾÎD�A}0y�������E}4g���hUt�o�%��vF�FIi�ۙ�l��X�#$�	o�i��\=�`�}�عū�̡�����Ǫ-�Q��=���ݞ��~�U��g�ѽ�|\�ڎ9H���WCL�����m1[�q0�yl�[��%��"�-�^_?��i���I���$N��?�f����則C�+e�P��(wAB�O���� .�8l��/5��~��T���B렍�\�mBK�.�J