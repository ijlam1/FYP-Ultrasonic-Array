��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su˸Y��'��d�Ay~�`�i���o3 1&����1\T�����	��!mF��
��\�ݘ�#X4|'�~a	N�1�""rϗ��?���ݝ��^��lt����d�k>O@�0�#/��B�#q�@�;<t��:�[-���&��5/(���{���i�9�о=�%}�~BW.p~+`�l�`��c�����eB0���iأ��䧽�|��b���f���	�%h5Z�\/M�`�i*iC�zĵ�0��;����(p�<a٣��9�/� ���Hǚ�Ӫe���5�4K�q*��D����%s�*W��;3�|�%��HI�t6�[�ZP��Y	�QR��-}�D��I=�.�,>V���R�C;�Y2�V)Ѝ�� �i��<����k��M����.c�j�ﵡ�u��¶�L8~���:`��֪:����:rV�ϝdB\8H�� �4������F�dٮ+f�sZ��t_E�g:�=�n�/���'#�EK4z�h�Fm;�{��eF>�_�D~&������t�3X�X����h�Ν�Ǵ�V�����+��ԁ][6]ӵi�Wۣ��2¬�J��.�c�u3h,�R�B��7J�/J�XZ/ʈj��p@�$��O5\5�6�����A�:9`�	�hL�΂�{��;R����.��*|�
D{����Y���]�6��K)�
k���ص���/��V��ѽ#�!
�;�$Ö����oOR�f����	N!TP�38kbD�x>]W'_��N1�A����M"Lg.$�U�jJ���_��w) �o�{D�8�5H����fm�;7F�l.Z>.���w��ke+\�2zaEaV�\�Ǿ�kn�o����Jd7�ӎ1H۵rT�c]�$�t)w�,raDQ�TE�uo�*��A��cjB��z��B�\M~\�:7�r�N��Z[܉��HhB^�?���í�
ME�"��f̳I>?�ΐs
I�����@���jLG�DFS�d���3�T[����,�U��|5?�P��6�8���t,D_ȶD{m�p?�V��&Z�g�f��}y�i"�o��d�Ya'?�*�	���r��D7j1���]7��5���/�t���A<��u�;�f������(�e@ŭ����Vt�ʰJ;�������Qg�4�u����|����6)�8�0k�e�P̅�h��ٚ��ӉS��c��ɷ(����1��΀���Dg��1���O��H��;D��2q���!�S��!X-u��� �힂Z8�Z���tk�pu��S��/Eh(R�����a@ѭ&6c�S,����͗���R]7��ˀ���b�*R��j�;�vm�x.�l��Hq�B�S���ͫ��\՝�%�S	4�3K�:���D<o ,��v����|�_����[$䚀f"��GO�+COj�K��2bUB�0����"̓1�!]~
ex���+;`����{�4,<Z�]o�H��t^6��%����Ce��G#��tac��_�pj���ew�U�+�#�����k	GU�{wtfmu���fC�#:�s"c�Qӡ�H�G��W:��j��3C����e�i��d��L2p:�b��hV� 2O�
G�uG�c�CW�j�)�@�IS��Rf�E���hq������%sӂ[�Qa�Y�����0������mh�|R/=M���d~S�V'���6 ���Cn�d�� Za:o'��K�y�fJ��S�7i���/�o�9W��)g6�I��Nb�::Ѭ�ֽܓ��.I$h�=�,
L�����1iQ���#0O���p�k�o4�AΚ>�H1�J�e���kaB4�!V.�&�;
@
;�Dv������XZ,Y`j����7�����`J�a�Y�,�TB�V&���A�d��B�������KliUUkyb���N$D�$���@����b�[[�\�핸 $v���2����N�z�k���]�n��{��=���q
@|�.�)��/����@ ʇ����߈i������%�6��6A����?ی�-o�#J݁å@�}���w��� \��,@{�H{'�zD�Z� �&:,/� ���ل�a��ğSc��20Sj���7�ݑ՜��3ڏ�(Wf(G�&塷/3a����!����Jk�X�$�R'���7X���P�f6a��\�7��z�웤u��B���mT[���-��W���ê�-�_�<6�,��u�"Z�����^�ܽ�%X '�2S��D�j^�
���Lm|�E����B�M
��7J����0���6c%O��M%�>�f�>�����m;�����r`Ï�	/�Һ��a�^�:�H�Yf�����@r��*�1��n�\:y/.����*�&���X�f����m_�˒�Ϳ \[�n�8V&�{��&�6���)"Rh�����y2�X�]a�	���|̣��P�3���د�+�K,N�z�N�uJ�H�e�v� ǧ�mu�p�������54��:��������ĥ�C*L�ޖ���u�BU��n"��Ǣ��D}��]��k��س�Q��`������X��QQ��*E��u}����fm�vq]A,~��*;��r�yC?�9?���DF�AS��猐����_��:v�0��*k8�;G%�����twΦC��
y��vç�o,�`ŤO7 fu����6��|�/�)�}�ڌ�����t�i4��˦Q�ZW^$��8K��g��N���_�r����[gn�a5wd�%�&��U�F{�Eqwj��S����v�{(�k�����SXݳ��,��FY�M��nz*�@ԳQ�n�ko�r��aG���i$��E�^.F�='&77����{()L�ej��j��A>/�EyWg4���?ί}�':u=�P()��P��>����M���Y�aԂw�i]	e���%~,��� [#W;b�K�0b���-�<���ݟn�U�:�A����^aw8!�n�X�t�M���C��c�T��DcQq��t���)�/�S��̽��v}�WO�z���P���-����G2�`g'�Af�X0W�9u&]�s����5}�g�5:�_g� �ω�\��UVsIXp\�)�BK�S��,ֽ`n