��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su˸Y��'��d�Ay~�`�i���o3 1&����1\T�����	��!mF��
��\�ݘ�#X4|'�~a	N�1�""rϗ��?���ݝ��^��lt����d�k>O@�0�#/�����"WYj����i� �N�7A!�@<e�]ң�;��5DXL�%�����f�"|���\y�]d4�V���(h��_Ϣqn���RL�/� 8�OK���a�Z����IL܅T?5
�Nx0��Ϳ�7͋)]��2�� ���S-��<�&42OƱ�%�N�H�s��)}��Lo,����;��?��'[\�W_ ���������=��hm@W�)�c[~+�!?�3�.�2ƟN�[�fx_�O��[����*W�0� ��������?�"H&�� W�y��W��}F�� >���hfO[A/.�b�N�����c)��l:�O+��t�'��k��OD����w��o2�
����y7���Z�!b�T���3&�ϕ�h!�j��/�3 <X�ƽ���YXMe3�I6��2r�\�]|i�(�1�O,��]$E�®�����fT�rT��H�-�����ч�3�1��O����0TGۙ
�n���<];H��GV2�d�������Q��^+M^	�����D��aB+�{1��r�M�����@�)�F�
p�K����>w�V}%7�ޕ�k��n��)f�qA����H�0[�SwtvX��]�ԟ#`�j)�u�r�F'��X�QKP���m�B��~�lƼ�9V�x�r�=��Q�v=vðٍsSΞK����rS{z�4/�$g%P8Ęp�;�9�5	./�^��չ '��O�/�ˁ�z���za4�0���ゐ�n֤wFV/��*�rS�3��
��	�Cc\+f��y�M?�A�.�%�JE(-
�FP=|pЃF�b@ձě�>=�w� s��/Ǫ�O������{=��A�T6�6!Ơ�D�[���OF�l}:e�⮶h��u鋯;8^ߢ�t�%���9?�_W�t�#p��r�s��ͅ/���3�/yȻ1h��Jd����*���T�ב��*a��g
*�4D��O}ăx�������E��'�HB�\_]t�!e��E�u�`9��vLm�^]Sɓ����Y�A��l�L�����u�}�|4�<ei�ȡ:lo��m`��Md_��[� �ROG��@5��~����)�q9�@U�` �0&�z5�#����O��(�E�I��I��`X��^��s�����[jn^����T�(�^�c����[���qu �@PKq��������ވ^�����I�����c�~�h �-���+\U��6�9cXӡUOg�*^�&U��б>yE����TJ��vt��0�u�
�~�`ݲ���3�a�v%hVYm,�	��VC�I܂����/�ia�	?�A���ͤ�����͙�-a˖��>z(�!�OJ��/�z�w�f0k�M���K��$�P��R�Y��Y���ME����a{"�G���$���E�6�d����0Tl.OS?o�������m��t�/�_o�w�Eij��Ƀ��7ѕ�MY�U-|^r���sz5�]/��ʔ}!6���h��=���/��&g?�GKa>�*J�R��������ѝ�M�Bؐ͊�����E�PLnZV��U�	ؚ��Z-?� 1Ӆ96,��y4<u��zn�⩧S�g��%�ʑA�l�G/��x����H�����iL�F�)&v�Nu�����\��R���^'Y۔NV�f&S��r5�K�=~�Y�~����5�Y�z�gt܃1e-��e�'g��%w3��Q͑���[��%�W�ף����![Z
,�6�z\z�^�cw��|�����$��~��v5/~}
k0/����Ѷ�I,Ȏ�^A��J��σ&m��8�m�W��Z�Sh�9y�핮B8��_�j�f4n�a�]ދ�(����n����ʝ_��d��2�(`@�'��9���Y/m���p����|���sE�m��Ju
Ίz6-g�p��FB�I����g�^�����o��2��B��:񅮀��"�����"���p%l��������|��l�f��z]7��Y�LYo�CXJ��S�]�ւ��O�̉ך��C&qs�cQl��9���l
'��`l�/
���r0���O��[�����U�G9�o����h*=�Wn住{��-B�+s	
NM$�V*�S;w�.����o �4�|�-�P�"��Q:�<����3Z���{B�zj@֎����9y!t�2� ����;���!HwR`�P�
��Yg���K��,�b�yq��I�;��<���y�];V%n�����f�osP�:�6��ْ�%vK�K)�����"�����M}Z�>���HV�M�;$R�V�r���93�EL�у�Vf1<�v6���2�ϕ�EA�NH��>2�x}����E 8 *�0Lns�߃bzr���Y��~�h�L�:#́:bf'����%%�2GA^��qPXh�;U\z���{�>�È���|l�߽$ɼ_ҫ!ƞ�}v�v��榌;㖓�{3Vs�5P�Wȉհ~����bso��)�i����gA^�f����co��~zh���`�������?�J4�Q����!�-��;V_3\�%.󧁯Sg�+4��e�$�xX�ueZI�M���	&�c;!���qEW��<,�Ͱ�d��.�O�ȇ��*G H;#�*�ׄF���rS��3���S!�u������sL�����P���ٹhS�����+�-3F�F�Z*R�i��ǡ������:�Nc-/|�4>�	Cd(���i4X��l� o��Ħ)�u�+��Iiqd�«*$_�N��Z�tHN��0����!�>��@�����)G�y�Xu�	������9��Z
>t0��L��Z��Í �[ĬH�~{�$y(M�&g��@��vw���DȐ�˕�̓ ����#�).�,E�|G�r�� 7u�ʵ$Ve�X�{q�6�I���YH
5�c�VNX.}F�T���W�#_�;"0�I8�O��B����o"�_9��@>��˙��7��ݞ�S?�d��&�N�1@<!B�S���W-�/ߠ^@B��Y'�{��w3�8��]�˩�R`>JE����/�-u��	���ގ֜��&�e͟�v0øJ���͇��p��F�j�QwUg	*Z�۳/K��Q�����,�ҽ���4 "���4=�t�2>{�i�a?3��5&]pJ�R�?�*M�!;ʆ>�#Te$�x?��C ���w���/�Сt����-��Ʒ���@� �d��)�7?�zz:H��I�*�$Y�3���n4����v����g�mg��O���O�f<^1�����1j.��$���UH\hc����+2XyFm�bü꣉�ЉAeVLOױ�{JO,G��¼/�[��.}2��r�N�����+��^�	�*P�����z�H���� ����k<{����k�
�qo�����"	�罓�D��5.��!��
� �M��\eN��M0����b��� �ɡe/�'R�-��d%�h�*X$_^כM������Q��}[���7̥�"Ur�j��NM/���
�@�A^��9����A�ڙlֻ��.*xv������CGaܶ7�#G�YC5�	oF0�l��܄�(j���T]�YOc)��(p!�#�?a��>7��HK;�
;�eч�-��خ�am�Pn�y
����Kw�(����e)I�@P�6��1D�߫x4��hiBWl%�]�y�|ǯ���g�3���z^�j<
�����7�L =�%	j���ұ�W�_ ��ef�'��9m�
��b���?���y��/gl�C��tvb�ob!�`韞���OT��ꞹ��G�F���w���� �I������\�x�ԁ_hp�TX5��h���%�{!~�c}�-�·��	����*��Sk���C�G���F[6��U�(�"����r�&&�^��&?�2����C���k4�k ���Sgj�0ē`�겘����
)Y�z����L�,%��ZØ���=Ig�&Ԧ����!��{�%�I ϬCi�K?�p�k��`��A�G�z��"�����������(,L�:���͊��?���\�qӴ�Y���.D�U���R/�ʉ��՟|�yWZ�[Y�u,?�F���Ց�7[