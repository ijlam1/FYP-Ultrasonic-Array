��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su˸Y��'��d�Ay~�`�i���o3 1&����1\T�����	��!mF��
��\�ݘ�#X4|'�~a	N�1�""rϗ��?���ݝ��^��lt����d�k>O@�0�#/���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ���7�dA=+Y�-k����c~��5���BmgKD>�Z��n�'f��\F�O-�q<��3��3Ʌ��:>�u{/�~
m�(D6;���eUi=)�'ܼw�Ӯį�m+I"����3�UL:�\�I��b��I.�.�#5��E��klL�~;�l2�41C�ѵ:�q��хA��Α�PB4D���{ �0�!A�m7?X����=�wc�[�/�~�1c��0X �*�p�3U�e��}�^*51��r�H6�ڵ)g�wwoP��Xm^��o�Q[�%I#4��h�!J�l���o�{�塁yy����8��v����H�Hʴ��e7``dU�.�N�ʔ"d�ܐ��μ�y��\�Jجl��u�DtsT�Ú���8Q���</����3����j�C]\q�{8�T�ZЈ�׀�l��5_�SlM�Nqц���(��'��Ǣ:cX�wB0��e���_�qW`:K�E��1}�=���p��ڒ)x�`O�}f%g"��oC�J��Ż:���܅ˉrے���
.([����ي������Ob~O�3��C'�+t�aX��4�\b�~g ���V[�D���^x:���c�ж�:f�s�i��Qw�ք�g'�6���2�<>�)�I�P�����Ӳ�/}��ɣ�N��U;}�Fl�!��EX�Y�P}ҽ@P�9@�(��jJB�DsO�>"t"�ڐY���4u�Z�B	��N�3k ��r�H�s�gS��J���	���l���=�úH�X-��U/%pY5���_r`�Uê#�s���^Ͻ"q�����5�03K���#A�}���g��v
��?�q��ŁO�չ���#l ��0����lP�?��J���G�H�wWoR^�Zi
PϽ!XR�X�8���`�)[LNz ��ǯDP�W���:�w��`Ʃ1�c��1�N]Xw��L\��!�:���w�~"����J�y�6AV���,���Wt�_�`�������.�/x���ci�?X�HY�~!�U!hQ���{o
�©�>XI�x�#ܳʆ�$�աgq ����ws��̯@N���X����;L�,��0E�T���ʼ��{{���Ħ!oF�ŝ� �/�j'������HX������ӫ�8��yZ%�EY���$�n<J(7����z�0���De�k�\Sȓa/��|��Q����V2�y�P���n#�L?���L��6{KQ@���0�p��C����q����r�eZ.�%=Ga����31R�Ցi��=�3�U��34KjȚP�UF��*f�i�v~�M�| ���~7;��Xl��=ʓZ��ڵ
7�Z��>X��|�02_��`.B��v2��^A�p���~�W�FN?�Ԅ�%R�H���IlḇQ�F�蒾��J޸B
�W�����z�*��j/6��|Ա�%;��%��ɲ�]�u�=�������%�T�a7M����V�Smу�+�7yb��õJus�2��V�-��;�;2�3�Eސ~����{-�|�F=����~�^uO�<��ɂ�V<�dH�ɒ4��u���c�#���$��C��|f��s
��b����0ƃ�,��2	l�z��E�w��{�V��w����㌋ڥ�Jr���>���X��/l�L�Z���t�K���r2z�ឰ9P-�*0��<Նga���=�@�\�V�K0ϊ���`�9�A�je[�&	�T�Y����4Lz�<n�P@=�"!�ԜO{�5F���+�r�w�޿;p��I��I���bԎo�k��<����V<�Gx�Nh�}ɫ�$u��/U(��A+C2U�Đx@�WPIȶ�r]� UY�c-�A��V}���ٹ��.�De}�kLd<P��g�R]�7�6�@�ql��������.��NRfNޛ1��~�~�寢�.�ZqOk3+������f���$I�d�
Pw�˨��h�V&�y�Cv9���,Ʀ��Ȗw�"g��|����N���~�n�<R�;����!����9�{�޾v�j��r�0{�Ѝ������%�ޠԛT�N��DEY48\魭u�'+贕�7
�<s�QMjd$��W�!c}�2��s��[�l��X~�"����D�]��al���_"F�y�]ū�w�t�|Yk�����4��X�����K�V��`����~N�=[dZ���.꥔-���	�M��0u|rl]M�/y'��,
�LA.I���d���lɩ؄c�)��ŁT�x�1m��t�t�&\�U�������S�X��� &���t��`��[�+t���?���0�dR��4��������p���+w+W�3o�#�S���y��oЏ���:��k'�{B!Ͷ/��<#�9��	.<
��}�V/���i�༞Up�,.�E^p����g`�
�|�P�*��u��{t�2R��3n�,�Z\3T����WIQqD������\2׽#Dy���J�R��$W1��|��X|'8����G�;�!g�hm�_�P��g�@�t����a�/,8��Ȫt��r�m!��dA��C�>�/z���t�D����h��%�K����A����i��t�#*�HП�4�Nk5�?����5�=�,�FJk�����X���K�U	J}��KY��X\T���?ʎ�⮨SH+�g]ܫ�� �H�W5�'j�(�6e!2�t�!��s�+'�b�珚�ܕP�#�*{��-�f��x��D��ܶ���|u�]@�����#ޔ؛]�t]xmaGÌ`��1Jgry��������S1�����B�p=�O)����h�k� ����cmX$��7!ې����A}&��'ٞ�� ~I/�7qs-ED�Ӥ C �k�s�� ~�@�V3A�BJؗvGe��7L���^B��x�0'�~�� ��K;���;���|��Z��q�	>%�ߦ��}p]o=9O3r=�Ts���m����p�� ]]S��"�J����X,1�Ae��^�CFQ��h�'|��o�M����;��C��I��r�F�3����ɔ��M�:�b�V,s�[zf�w/�a!�P���N�ejP$[����#5 1SF��}?s \M��)�&͵3��h
�jY�����IlS4�aoR�S	�]�ö��۲4I_��9Xc#�=�Ø����&
_��/�9G�W&���`�~�HQ�\u���I��S��E>����@F��G�����@[đߑ�$g��4�E�x�)�����U�4�>K�ax( ��z�{7��9�Y�r�Lrgu @�p����ߔ��m�J�"!)����?V�uJ�$;���}O�b�=�ܶ�<���Ӿ#�-aQ�mV9�9���O�e~)��Cl�i��N��tscI_a�Ec��P��ʁ: ��.��d��^�=^h�	X�mGv����	@s���_�.�(��r׃�r��!!ݕFA_��
Y�M��������?�bvK��..��	�$N�4d��w��Z=�ݼ�:{&סu?��끖B�X��?�q�*F�>��e�ػ��_�_�ӭ�y"�5'�zF}#�7���)�\�8ػ|�ԋ4JŮFE��3�S �<�f;-�6NGY���b�����H/�!ه�'���}B�"�&Tr�c��헉)�+6���,��"?	r(UL@U��x�6Ax�:>8v+`~�J�}�E�/e�c=��ޗ%������c�u�k)�?�=Zc <7o�>���ζ�IN2NL�*�ٌp���02fL`�~�4����6/:-&�4�q>OƉF���z�󓾄?��3�&"}�����[NPd�|Ϙ�u��D]vi���^ب�ZD�ڇ�6�o�5[�?c!�� �U�"ly%�YG�$�!��R��AY ��b%�1L����KыG9�l�L	��q�C�K>M��Q^��
���}6������Z5������Ї��;У;1~�#=|R���K|rb�=��$��U��7��$���݌0:��dO~���w�TC���z5Wɣ���JQ֟[t�~57��!���&�_A�,#��o��]v�`��hHW��;1�^�6?3z�����@
v�S��pL�L-��l��s�l�"�}�ѲcU�`@�`q�.���[���5�X�� �3�+�Y��[2���<7Q+�� �6Wqi)%�xӁ1Jj�_��	gM�d���r�y��m��C�˚I�K��db�/wbx�B2�¯�$����mO�~��LD����h� ���g!�p�rj��خM�>[�R<"X_+�k����q���&>�d&2G�p;$R���B�hϓ�l��&cS�خ���U�whQ�d������o�M��ҩ��=>�$㗺�O�Z��N��:���K-�4�b{�Lw�9Ĺo���U�����v���OI^q$xF(�	,�9l"�r�'�\ì	M��7�E�z~�vp�N�.�	�;��U�R����k'�Kn�=�L+�v�	+rHzs�<�`�|�q'�&�{��a�ٞ�����#���K����+�G���ւ�ʜ������̹��W�<Σ��]����{]��ǚ��=K[���2���o�B�<�P�ؘ�q�_u^���f�Q��g�{y-��-�|U�@!<x=1���H�cF��K-沢�C��#��	t�`�>�r4e�I%�*kD|h����?'"��2�O	���y����/H	����kʯ��oh,+�Y���Ң,��e�5>�缝3j���Qȱ�i�!��\*y��>�-'c��e��ҕ��(�|���%���r+!FL��z�w�	t��GD��N�wM����j�V'�u7' q$�8_�EU��A�;O��<�/w�����,��*Y��H�Y`@yOg�5���}?��ܱ�t��W����q��A7�rl��&V-���ac�$�嘰^�����.Ok]�B��g,1��ʚV
���ފ=��.��nI�[�)��Ns�Q:��r�%U�0�_��J����ji3T�lA��kkgbg"�3�TAjA-X��A2�se��v�E����P�7v������њQK8�O�] ���0�W�]ߖ�N�X
�����g���c�/@�HO홡�u8v���T9�֚Ty9���v���oq`'Qk(N/�9r�Vu����y��K��YQ�I�<�CC���&?!�A-��qwO��/�4�R3�,68����_���uU��d���ck37q}!�8�Y�,o�����X4>YK���)�H]089yD:H�Հ;�[���;�, X��oU����e�ݮ��i��]"�z�p9\K�7�#:�YH6��ɴ�w���)��!5czz�}��z)��΢�̈́��)IV�0ڹN��9.	��{bN�\�`��2����d����
]�j¯�N��+]��Y�l!^��cQx��7-��j"9��1���
�+2���&��Kp^�����w���O�y�r�P��ҲWtO�|��h���C+YL�hh��Ӭ`)%CB��	�_�W��Dﭣ��7+u�&ښB_+�Ak��0H1Σ���3:�����,��K:'$�k{ۀ3Pi�x�ޮ��(w�j8�sd�C3	����[FX���:�EJ���Mg;�[�o�������L��Z*��ϸ֏�<ơ�W�A�sl����~{@	!u�kk��2�@�/�F���	�M����@u����4-&��[��@�Lj�-�m.hK�#��@��.*�p�{���	��d�d��?7<suk�a�{-c����#E�J�<s��RV'�����2����(�p������/�<)1(MO�Ƌ�!/�'ӽo&�;�|�A	����A!����K�O���)mYT&H�x��cs[�=+t��Z���M/�y�ahIx6���_7�I)Y��*Pw�nH@J&#m���Hv���jU�Q>����>���v(p��W�m�e~2|�qԺ�(gd�bD8`�e|���z�c�n�ZDs�ؤ�%X�| I��6� LZ�R��]9rw�DsZ����͕�n��������붟v)�̟�o��jY��0�@@m�����i7�E$,r_cy���~lc�c�Ď�5sB��x[�J:��X�=�����!<V_�D�ZD��+t��T��m��>g�H�[.���Џ���AbB���O�!R@��\��e�F�+�%�����$3�i��U�$�t�F�����I�A�'���h]�:'#����y��5���6W̖vwl�1T�IW�7�B���x>�9��� ᩷8M~��?����:��a^Qe!��&�,���W1<��rbh�o�#{�)�fV���>a�Mw�n�c��Ѿ������R�����RT����XF�I	1<��G����!�Y�:�o�J
Zߘ-R.~+�@n!�%YcU��-��uDP]u�Zl�(��2 �k�>+m}�=�*-����9/�1��h��?yv!h����.j�3�Xfe�8�����}�yN���:/mP���� nJ>Õ02Uϖռ��[J��-Bj��T�>� ��k������Z��
n��C	�������l�-�u#�������g'>�~3���|�� �3F�� ��v���xE�����*���������G	�[ba��h�*0���r������c���>+��
^錜sx�cqse� }΂;��4�4`S�7,/f���8aW����>!��.*J���:,D$�؞H��{�`�o�U�w�0:�>ȭi�7�_/AnL���"2�+L/r�"��}�/��iԳH��'4,`*[�D���A��8�S��U���g�Y����b�oF���`7��"��pc``^��IK mv�)�Pm�P�� p݊&u�bV�	g��u��������fr��>cٶWc��nF�.����?��n',�XC��v��מJ�2R�[�	p�խ����X���<�k״���m�09[u!��_�9�tIV6�i�x��ɮ�T��Hmrd�ԩ�{y�áiQ2��4}�0�4�j����	���k��Q���OH/����S[ �|(����A�o�'�q�����h$���؃�0�F��5�{��Y~���8��I���/�=(�YP�����؊�3�E��0oGVY����|a1w��YG��fT����Z����r��E�05d��艑b��v����+;�5��*�j��G����r<�h���C ��L�@�9�q�FD8j�\�C�@/k
Hp�w���k,��S�,�|�>Ps�����[�ˊ��>�6|���}�oa��#Eˋ�:,�z��Z��E���� ���P�ɦ�~�ϣ�.�G��>����v4/(�qMlК���dnڹ�� (Z0�E(l��>�|u��Z�4��g�ӑF}��t������?�����qkz�����9�6�3����`��?����3�; %��L���0 ݷ�K�=�=��A"N�Ĥw�<֜qr�vĐ���z��A�^��S�F�H����M��\4�e� pF���­/5�լ�D!A�5�1S0�����]Ar��ݡ��;4!��~�4n����- ŉ�릏s8:#bvu��V��|��u���&c��+ۏ=-�s��B�㖱���:�M�+8�B�� �X�'Vi�,�y�=R5$0����k1�(��ݜ���詇c<H0�M�jw�j�"����\q��
����S9&&���iO{=��3@�<ɹ}i�`��1ñ6ɰ:�x^#�������.�Ͻ��,��.H����i!"���� ��^m4���ʸ7�M%S( *pqD�wMѪ��x�$n��BC�:�W�b}�cMAv�I�xio�O�n�r��Y��wxL�Μ��&�ֶ	����l����8c�20�G�h�A��GՃ	���K�Bє�������q��ءZ!�
���'T($���_����S=��di�d�ȿL�;�;�{�Xu���fyE�������>S|u��4�\Z�	{����/>6V�ꊲ�f0E�yl9�&t�����I��}��,fKEn2��V��"OZ���}]��"��U	lԭ�g��Ƀl��g>^�}t��i���+��������ٳ<a��_�ZޜB�
��,㖼,eSk��b�D�2g=��Y�����BQ\�;߇{A\���.̺ҥb�'����!��q�c��ϟ��_��
^)b��N`7#g`n���mC]�$\����&�}O4�!w���Ll���!6��L�I���@�$�Fz��GaT�"'z_O ��}�)�����u��ڥe':$�����*��${�XT�6/����!��l��Q�M��t��M��߹�Ai�P��r���G���搃��/�zǸB�}�b�`��´���'��b�p�>�,?%�C���*��	[�ߦ�x�P��m�"�`��c�3!��%�<�[��(S	�?�ޒI�KN9*[[ܘ��MV]�0b�2$n��/�s~�.����0�K?��_P=��V������TI�">Z��`���	�2�
��<�򒳵���g�mlAG�غ��s�/~K&:NCfY��g�y��Mm����*h�_���FÎG ��nn�&m�i�;c6R��4p�ׅ��T]�s	��%��?��US�R�j�l�an����|���
Lѣl���F;��O���r�"I�Q���c��4h��v(ZO���	�*�K�������[b�+c�:�'������N8�=��1Po;��s��!@�m]FR��)pu�U���Ǽ�P��3"�5��� �	�Ό�ϟ�|'�0'�2P�Y)W R�k�L>��"٨�\E ����ߖ��u�qX�Owfl��˯�p�o%�=b�G��n%�/���C0�@v��{��)Ȗ���cT�'H���Z�A�:���A��d)��pP��!V�*��$�E�����J�1VG��Rp�ud�	&2*���z;�0��*��#����;k��x����$��uze:K��.����ȁ�3�4��U�.��x��%H� ��r�l	D���Ɖ .���[:1��&��]7�<�3R�}M//A�'�!Y8���}�~�N- �r��1�g�&Њ ���S_�sO�>O��sd�q]��]����k�@98�fVks����Dr9�r�̆_I��G��k,�Q���	r9�M&�M�>ܷw?)"uv.�z�b�W���p�O9_A�k6C\ V�� %��a�O��I�+�5p�gc�S�!���--9\�|��������uc�%��D�S�F=�pN
O��_cըh�V�s7����r�9(�̾7����ƳD5��@y/,�����23�q��O��SI\p�����!}�%o�Ñ4T���PT6sY��a��F4Xeu�-���� F7]��	=Ud;O��4�9Zq�{��I)�0���4kȎ�>�����`�A��=��=��&�p1���(��Q�[Aдx2�������Pk�ΪTq��w>:���0��1�Ӧ� ܌R�T\8�j���oM���A��	n3u#4P��6�����f?�rO�#��#/��Î����\��"�S��em�����y�%Q��[*]~�dc�bX<j��/[oT\���Z�-�A���LPJ�Q��OgH���ek��|��?���W��67�����u���,*��r�T;���fAl��纴��)=%���.��&����x$�Y���۾��9D���������w۱G�HS��@�R���*�ȓ���[̓���� y�+�ͦ�F�#@4�)HXr�;��W���Ίf�V���R����W��_w&i�md�-���|����2����r���25m��f����u����bF@4F���l"�A�i)iM��q�7��QUM��ޔ(�i��)�Bһ<LVE�6y�l�7!JJ);��|dy��T�kN�����ǖŶ����b�L�,՝9a�B���}s��j��k�������Gm�=�x��-���t���])�k3��f���Ň��ݣ�h���+)[5��t�#���1a�C��.�Z+;�͍v��+������r�"A��vO,JZY�+f
�h{j|5=�<��p���1 uKZ��� �v�Q�xQ&�{l�6���ȷ�jً*3Egh�$��K�7nL%�v[�5��@%���6q`� ˈ9?{W�,7�P�*i�0�Q���$?�a��O5�>q�ed�vH1�r�SU��0e����H�Ű9�*5
O�Fw��!:B_�/ڌ�p�r[�'|w�S���~�qh�9�zˌ�J,$[<�1N�͟��o�B0!<=W���"�/��=��D���"�W��qp�!6:`�6��������>�;��%7���	�y���k���4.sQ�66?���^�p��Y����Z6~͐r۸xu�QS�&�c�&j}J+�����<�=�ᓗ�Ov�㟧/@4e�	ə:�[��(W���d7y"���������q�u�~^��L94T�8�꧛�̸8�H	̹�'�Th�X����P��F���9�����d<k%f���uv�o�9{�TE�a0��RR������+-ۥ����;a���#� oT*i����Z��1X��j�?q�ѫc����%����;m&��Ϫ�;��IR���SP��2Kp�`S��ag�hL�����gW鈭݇,����;8Е������ө��D�������5�?����"�?>pp;���s�YZ-w����b��R���;�n�1\���ֵ"KmJU#Q*X�\�9$�h]}XG�x7�Ƒ��*$��|�?-=�J寏�.�KP)��^΀�*^֯%<csA3��;`�՚uD�8��d�U d�=qY�	��vˁ1B�h���vw&��fY�7�u�(��G��!���c5�F��RfO7�E6���{�\O`z9���zQJk���!ez�J����J\�H�軮���S�Pf8�i�(��,��1���Q��Z��I����B9L4^0n�y��M ��P3�\���RI5��]:A�VM���U%2d������naH{�Y�]`����!n�]U���V��0%�MQFF0���>���b�Ć	EGTJ�K�qx¯E+gW����lkڟ.b�������{j�t����"���g���˴�,?�o�>�