��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su˸Y��'��d�Ay~�`�i���o3 1&����1\T�����	��!mF��
��\�ݘ�#X4|'�~a	N�1�""rϗ��?���ݝ��^��lt����d�k>O@�0�#/���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>	��։�������7�{�ߑ��!#���
����8�[h���}��,���4T¨9��8wU_���a���el���`�//��&Q4-���j�竔���#��G�V��"��~N���V:x�
=~�	��9=��R%��V@��a].�<�����B��v"]�e��:� �Z]6� �ֹ(��gJ���������'⬞/�tO�"��''��P�\���>��pi"��/��b�������� -N�.8�[b�#��H�U{��|�ز*����)-d�A ��.l����*�"6;/H�eD�w��X��ɮ.kj���
8�ŋ6�b�A^b��9dտ�PK<���9�|<�)�]q��8��`� �g�ԁ�T��_�Dn6��o"1���r.C5������ѻ�LF��~Z�ݍ���˪Js^��>6V9�І{��Fʋ�����n"jI{�Υ3����`�R����]��h����H}�vD�� ���J�B�^Tk��G�ŕ�C2 ��GY!�n�#�d�4��Ж���u&W��B�`�B�1��Qa��Al�fNL��s)i�a�zFIT$�6EH���LHD��X}�2�U�M�I�Tc�?�yK:ͥ���L��8�J�$.�I��Z#�FpY���K.}:��Qpb�F���J	AyY`-Sft�n@z�����G�ܐ��-��n��*��䣮`�jKNhf��k@-�{�|�����|jC@�v��غf�
�����<��H~�^�ڌ�e_T�r��F��iɅL&蔭+����0A��2%q���vT"�Sυ����a�#����/R��7:X��8_ћ!�>R�o�6�%��gcsN5T�y���32b����g1�)=p�cc�<�P3��J�E#Y�������ֈ�_q�\Ϛ��)3ϝL�vq`�����E��7�UC(�a���QWcN�n���O!=��J_r�iB�	.�rޓ��~�����'#�~�N����Gސ�u�=�Pvgs�X�G�\]�Yd���j�C�t���J�8��|z�SA} G\D��~(Vǚ,��s��8�P�[�Aeh�P�b��$e�����2�,��7�a�*�ߧ���f��h"p�Z��2���\2�P�����7ge��F6o� ̇n���)ג�����$���ò��e�W����p�pƸ�?�f?*qU^��忠࿻E�Z1`�Y֑�Y����i�ۑ̊'Js+�x�To=W�,�`v�+�1k�є}�^�,~&U%,�r��l�-�zꞰ_�uX[b��Y�Ų�44�{5�������J9�����l6�7��鳄���7'C��%}�%��,*Z���`�bx~�׮^R��>
�n���%hWH���7���fi�Ԣ�_�a����]��{����	0X���gܳ*^-}òPm����_��_t���}ޔwG^�,���x���|�B��O��~	IS�9G�u�!��'bɼ��9�Z��������
��dz�M�x{��O�+���s��#�Y^������H�>���i�Ã�R�I!"Z*x�>D~��R���� p����X=_�|O����PM5�����z���$�8���r^F9o����Y�NBy���G#hɥ͵#�U�H6v��agtȃ�tr�ɹ�9�(����#�;I���P�6�7�^o��
iCK]"D���8x���J����D���_�U~xa�r���%K�.��m�ܫ�C�� �n�lb'T V\�������
����9|��c���M$�Z�1��eD�w�+�W�Vw 5�'+�KG�~]
}�T~���ާ��J��h�7
LJ�6|�j�闻��)�3��ʧ���{�k����� S�Qz��B��-+˫���G]*�A�%���#q� �K�t�Nf��
����}w�547���]6�}
T��1�� eHĨ�Bf� B-�9W��=I<ȫj6J���`/N���Jy�&z��+L�ZV!f��#ʰk5�R���w��"��׿���+�b�	r�E��:��Z�R���8�\l�G@g_TXȉdx�CI%��5B$�q����|�wޔ���k@X�ϝb��p�ӱ�*kEFbU����Z��Ђ:�ތ�N����Ma�h�CD��+.2�R��4�狯�#���o���B���E�e9�`4?C�Y�H��%'t�&Wz��~p	�N�{%�f+�����6�K�����R_�Vm*�X��0�V`�Y[�i�Iu�o�\����7e屘���s8������?m�������6��Q��|s$�s�M��I��W�MLW��������A���G+#��Is9�BM
fU1��[3��?��q��響0�+x���X5!'�F捃KmoW&�o6D�v�4�g�j�-��E{��+�ij�9�?�K*J\���i��c��Cȝ�s��(�V�4�g�2��9�	����v��5��Q�%)�it����H3�3K�Y�0h.�V�"#K�{i=Q��N�U|�0����^��I�T7Ҧ�G�֭��Y��W]O��%B�`�<����B��J���pZ��x竺B�ߵt�3���*�_L���xṗ'��r��J&�[u�W[_B�,�	�)DT_d��]��L��v49~|��D7:�r�ɮ��?'ϝ�eo��yjS�����J=@f��xJQ� ��$�ν��d��h������,+62yJSy1��P�@�J�ޜ�i��~Э�o���)4�j���W�^�旦I|�7ɤO���Q�x>�9Ɗ�zG$����.�*�v�Na�yH�W<Ip�Tϲ���,:(ԩ��gv�T�zaol�S-[r�
����~x��F����q���; �	Ι!K�Z.A�2
�3r���8���ʧ�$���FRkpS� >[��/�^L5�4<�h�{Sߵ��.��������h�Y
~GP���2�k�4�Ӕ�/d��mq�ht�]�k�Hn��)���֐,�
�̆H�恘���3��ٽ	�?��x�� �#sj��@PbLJ~G!G�"��A��2��jU��S��LVPf���}y�������bz)֙�4p��_�O�Q�BbCK���2�X���d,efw.=��"��T��UYa�3"���X`]2v�($9��rI43y�����U��X�LҀ0.�d�A!��'o�<�&�����O0�mmQ$<&S�*�_������}�!�]�����%2�	 �j���V��ˠ]8|[�l��TY[��R�ow߃��c؃Z=��?��!�<Io!D������K>�<rhPTEHv�lcϡ�������JM�"�^vd�Bt��!rj�	�2�%4��i�:6b`�YV�j��z��:Q]Gcɴ�s�_���a�a�tt��������[��Cņ�B�9�]��Ĥ+J^�N�l'��>M�Lk������q�=m��g	&�η����P�����e��1���|�B.��F�6.�n)�x�zg>�PWp�&g~a��e�� �>c���H�0q[���`ܣ�G�Te}�î7���z��&��oc��	ж}��ŋllk�)��}r�6���
'?&Z��M%o�l��@E��d'
m�����n��k��
3�S\9������몽�G�7��ޠ�E�0�w���%n��Z���˱����1l��)ˍ̴4�j�'��G+�	�U�U*rپ���i��i�v]$�F��c��58t���XG�L-�yT�����f�svh��7��Z��G%�
P2KǊ�V<����#<�Q�a!��ҟ��G?����3�/Ɩ&Z�8����9H�	��#Vw��̈�z��є,yF^���qz<^]��ut�w�C��	���������^�c��;v��0�ŵOK2�X�i��emcE�`7�����C�!����n��'6\�������!]k���.�*Aט��il�N J��8�Uӆ��\
H�:�������V{x8lF�R��2�/���k����5h�ЗOF�������Z@"�w�L�E7�YAw��+���M#�F���}��TT�LҒ�*F.Zg+f�bC�W��k�D	|�	�~�/�z����j`�8�eP6nS���H\���H��|�}'� ���bЁq��K���܆ObQ�j�	����O�ֲ���>x�g�􄍒�a�oqx!�÷���v���ȕ����o{���u���\�SaQi哬O4����ƏnI�4���AU�� ����ca����$�j���ܘ;�b3hz�*��b�	��]�%(��0<D� �1(�\�;9s�t6N�_&8L�J��?(�d�IrJ�k�hY�`[	En0g�7V���x�j�K����n*���\�쯝�m��K7�1"uK��\�"t��;�bK9۬�˭)�ƃ����qO~]���z��Ֆ�,�A>!C{P��E�6c��P�B(�0�s`��0��$�]��E����X�����
?�~ɒ,�J� 	
�L�nNp�{�����O*�HܝȚQ��]G/���*�v<�+[nq<��,-��2�y;��Z��1-�b�m5D����z0A-�����o�S@�K�ƚ )�4���wj[	HԎ�w=��h��eY��u��dT�&��u|0�q�Ɛ��7�*t	�b��w�WՊ�h)}\����3�>�|��<��Bg���b���l��Z��0��y�in7����a'��3����}޼o�zP�.1���~�~���V�gD�y�� E�C��u�Xdj�śc�T���f��9�m�ma>P��ɒ9����Iҡ6茉�%	���
z�����b!x\2a��*QfP.G���z���=��,tM;E#^�ɺ�ƻ>5����n7G�8,m���_�3nY�(|�B�7�i5��#��3�"�	L��؈��v֮�vw��e�#\��-�[
�)�0��g����-�%��﹔�8�O��噳�ӡZ��EU]`��7��ep rP�s@�.}~�h�v��HU���¹���.���Y��1k��Й��*�m������ð�U��N����^Ɛ�����Ŀ�t2���҂�q4���<�$�Z�Gt,�k��4�<��n�'��ϰ�����!5�ϝ��:B ���E�&��3���S���;(��P�@�����K=���A���{2�
:���mF̨��g�� �}G�bE�x4�ta]f`i&=7vy�6cD��\C�Da�9�-2�&��l�W;�$')�	�I�ň����
`��ߍ-������R���p�ܢ��,�)���B���� ���nkR4��zU��%��w(�	��_p�`���D�P�C��;�ί���i���u�Պ,86LckB�:8�ղ�y��Ԅ��]Q)OH��i�e� Y;n1�Á�yY�lq��i�C�p�5�G?�ℛw�8V��~����i�e����b��������YBN���""�&���7�mh9�5��{�i,������f����*����6�Mӵ�)��S{ �x�;�{m��'}�i�� vJw�;��4���~��e���Y��G:L8�I_�+%�ol�������#����V�Q��'i�-*6�5��CC��`Rܳز�B�|���5S�'�I��::���B��8���!�C>_T��}��qh3�����O������j�Ѭ��l��g����#ie���qVf]�t/�(���C=~����	P~//O)CH=<��@��Msw͗��M#��z�D�n]}~�%г:�_�R���[Ͻ�O�����70����&��"t4:�e����G�*�i��×��	�qt��Hc_���UTƒP�æ�+mA����ԣ����#���?(�_���O��3C
�Qa�.�D�
�(?C�<A�ª���_M�|l�R��	�����q�o&��NY��JBSC�e,n������ɝ�o��" �͞R����;�yY��D��	7Ukw=�z�����Z�tW�j���Q�^ظ����g�N"E.(W����������Ҙ���r��\*�TFη$�V Zc�b�_Y�`����Y�BO�{�ە'ȉ�N6]Y�0�4.�O�H ���!�`Z^{�������S�������,�*�O�e>0=�Y��	�o��i�[���ͅ��ኇ��P�����ҍ�����՚��i�,Ʉ�Az"�\lQہ� ف&��c�����]D�����R����z9�k,��n	�k��8��5B!5�p��XMⱮ�P$�t��J���?b�B/,���^B=!����b�M�ژ���]0��A#M|��*_�hy)�L\䞧z7�Z��_�I��e�w	��m�]2����S78N��/m��u�r�(R�����K�7��
�&�;<G8�:k��ޑ903M�RL!�w̯�t��9��x���dâŇ|�lq�lNM����I��j�I�R7s�ͪQ��-
x���������cyH���x��d��(6���,861{cO[�E6TX��+5eZ=�(0Uy���m��ŗ��R��Ϧ%��
y���5���V�6e�;q��~=!�l����GT��6A&���1�5�}=�g�������H2������>�2��ؑK��t�fM9\��W��N.���t��� &Xe�1�s�GE�&�cdm.����PY�������Kw����'�[ؔs�XpK�l�[4��
�Ve�|�����.�J�W~����Ұx�']w�u�~X�r�{Ex;�<M(��Z�=��x�l:�NO&o4E{�g�P��.r+�N������i��o�u�~r�n��(	�3��ٽjYJ��K_���z�h��� ��W�9&ۜ=)޳?/�U�����2�pâ0��r��^z�� Nw��i�9��(JsJd�s<ڏ���}���Bm�$Q�&P﹌`����e�E�{�Ǭr����`Jci)�Q���k�f=D��8�7�ܦC��'*z��x�\�(fj(6�UP��N�ͩ�0�j-Z�TBW.�t���̷���2�WV<m��7��(D���)b��M���1��Tj������}2E�Ɂ9����AN�	ȡ��+B.��ټ#��(�d:�*D��E���k%�>�H��_|*n�f��OB>�`����!��W����y
Ě�����^{l���M�}{�=�H�zz[}�n\]n������iخ�H*�C�x"��o�t�Ǿ��&�X