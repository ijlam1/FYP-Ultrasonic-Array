��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su˸Y��'��d�Ay~�`�i���o3 1&����1\T�����	��!mF��
��\�ݘ�#X4|'�~a	N�1�""rϗ��?���ݝ��^��lt����d�k>O@�0�#/���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
N�m�H2
��j�Y�? ]r��j�p�V�d�����띜�7���{o|��hg�EbVS����K(�k|@g���)��i���7�b���&nDo�/7���)�&	!%�Kw���qi����N�c����S��g\<�e(͕-�T�d�G�KD��P�j;��|#r����l�|�ݾ�SQ�w�v���|d��2�ښ����g�Ti:f�G�Ǐv��3O�o�d��*J=�#��IX\�T������2)�En���3h,8�Cg�-T���9�αI�4;k���N�� T�"u���P�aT3��4���F��x��r�gav�m� �ᡟϴ�^u)].i[ݤ���*�X{���db�#h�ϟ�j���(&>����,���1=�<�-�����ơ/2A�_ o½���Egi͡8�Ss/�S���5p��A�H��)�U� �aI�Y���C��u�Z��j��-��19���r��WbJV�������1��h
W:��u�a-г���D^p�V���l�U�n~h���ĩX�ӿ�o|�� �J]�d_O��V���G�>�!v�}��b*����?P_먔o��e���a=�d�C�r��&u�'m'�Vi!21��h��|~���Gk{l�?h{ۀ���*`X��E���q\� l���)� ;��c���߷(��q
�cl2"f�t������'�ɒ���+�3��;�����-���2���a��4S^�w�)rm����>�C��(�O�nV����ww���͕��ˀ+�WqT��
P�6FT	��V�����5����	�wK�9/��'��_��?_ra\d�ll<s�5��8�ɳ�4.	�PO[u����z$���F-�����ٝ�eBc�g1�=�E/��i�Q����asO�=w�׻�.F��F�^k�pk� �ք�?'�v��K_\n'b�u 4�G�oגџ��J�����\^\����F֕��iJ��͜6�Ҭ��0��EІ%$m8��3�o�����[/O,S�D���
�z
$��#���sK%�\���7y� �
ڽ�u[�V�<0�؎�Y�W��N�����9�d�̳��t [W�����
�3�K��Ð��� �Iތ0�F�xs�γ��u�?2�{؄���Ě9(�D"��i���3^�y\�H֣˳�'�I��h]��=���S+TBM�al�m��BR��8(t�	uM�4mYڶ%����I�@��hG�ϣ˩qG��邼U3�X�lp)�E��l7}es?��U�%(!Ϋ!������{C�z^�s)9�"P ��:�"��aH�ڶ0�R�e�c�mP�P�� g�'wt�u�6]�
��ԒZNӅ$bĥbe��I�A�Sʆ0�w݅'t�C�L�ِZZ.�l5���]�ؑ;�uB�z߽"@fE�*V%��dc)T� �*��fj����)�I��o�Q�W��+�^4؋%����*��Yo`�ﱀ��t��a�nΑ`�r�@���b	w��Y��j�d��C�D,��EH�| �U�Ѩ��SI_tIe�-�K�.<^}�]�>$�W��oK��(�Ώ��:�Pi煒p4w� ��ey���^��|H�L8a�v=�Б�[�a)���*��<�:J���9_>Z,���f�D�>�]yeuf�΂k����7'���TQl�
�=^�.#�l)H�4�CK��0�� �c� @���hEG2��p{%��E�U����Qw$&Y25�~��CsU0������Ӏ�SɃ&SL��E֔��ff�R ��q��9VEzn�z���B���{i��C`�$�����t�I���`�ȝn�T���+����>K��z߻=zHzޑr�h��q��T��/�wf���Я��}`;�(��#TZT��{���������<��*��fXs�j�����V�ގ�J�"���XK0�s��zB����od�i��U��i����g�H��4П@Ll>@��$����.B�W� ��R��{�dܕ�Z"�`l:�si��j�,L��2�5�^��eҿ�ӽ4)')���G�HO5L��F/�ѓ=vA�N�xM����8C�������@�xa���$�m3�R�x�z���m�����US%��u�;��z}|����dОYÙ����y��kD5o��
�Æ]5F	��Ϊ7�0��bd��#�NHC�w��B��r�l} l�o��מT�,���D�$�3�d[1��(�	OST�y�jBY���ơ���4��f�?7���v�"�6c,������ ���R�#B���;��������ٓ�-T$A\)Ց��v�0 �i����jA"�������/���D��o�α�E@6�S�SM0?��u?ir��)}��#Gd�Ė�,�a�}�eQ�����s\��q~�o�ܑ�N�z��|7�^�2�먣�Cj�~O6Έ�
G�;ٸ����U>Ic|�i�8Ź���#ئl2����:ׯ����1��mE ��������$}�%-;ߤI��,�����|a�2w֦�z�^`���߬�F𽝾�����|. ���<�Q��
*E�2���G���Ox�u�n�ye��ɰp�4[$�a��ֺf�v8��@y���pf\���%��#r`+U/����aG��3W�j1�_W;#�f1H�"<��� S��XG����~5��,�=ڨ�.�k e̫l�����;�Q=<+����䣖΋=<�������$/�]cD6Z��s2=��-ZԠ�ۗ��kh��Wr@_f~A1FM��
 .�J�9ߵ�+ֶ͟{5zo��9$����'��ëf����Â�R�Iy "�Y�{��&'��j��_m��3e�R5����M��e���z��.^�v�ye1��F���g��:��A;��=I:d�尠2y�G8��͵�� ��!/l��L���u�y8J"L�M�F�SŤ����o���@F;��g��?��OL�tu~��"�&b�Hf��]��L;./��;nDf�x=�J�Y5�ֶ�`>nT>2M�?6O�7�J�\���?IK7Us��#?�K g:�2��F}�4�<j�>m�<��\���c�O�Xk��A���򐉭q�H�9q�Qx�" ��ĵ�"i�J6��P�MK�NI�Yұ#:�L���!"K���1�2P�R��#U�,a�.Ok������w_:H#��u�Uq����u����V~2�g�Rв�C<���4}��u���Jte�S��|�Ҋz&�<-����@�7�`�~1������.�9��3s�+���N��L0��mH�n@9!�e;a7�t�[�m9��.�懭�\AU:��r�b��i��1R�q �I��ǀ�����Y�>��eO��"��(��q��X�䞆����5K�8���T��Zr���d!
i��F��|)�wQ�FOR��p5`��\��sԧ���Y��S��Եq��ۢ]��E�_��b�8����Yfq7$g̵0l��i]Y�~���#�r��2�N_&���W>(F�`�k��o�W=罠
Lc�����L�b�3K���f���\�0Q^M�1w(�� b�P
��D����!��O��Z�|�%��Et#�b���
Υ�r�ۜ"o���^��C�1����h�7D��ga��H��-�O�Y�Z ��,�:$�:mG�l+�D��![,�2��|z,���&���e$EIp�����3|�̶��v�����"�2���u$Q�h�n	.ի?6O �x(�����n����Nh�;�2���
�=����-În
��K y���i2WA`bi�Un�
I�3��/;��d;qt�˛�[E?m1�����ݻ��� f�|(j灞�Z��<�mJ�)Kz�Ks��U@�y�U��a��m�gŸ��<��o&�;Pܩ�z�h=�����	z��_6���\����&w��
k�9d0�X\7<�)ؙ潢���e���N�<�G'?`�5p A�l�F�f:�`3!�1�z��Z���e��k-pq�:�Md���S���*	��Tc� XQ�傭0ۘ�RPI~�j�q~�zO�ˡ�W5]���[�RJ��&�1a���?��9�k��`3��]l��N��R�����g���ܙ��[��9��8fh@[�w�z�8z�#�f1uh2S������6&(7`Z�t�9�ٙ�Ż&�^��GqSuп�?�'�hW��h�@*/��@�<s�cJ�n�������<0�_t�4S�5�Ȃ\;�h�9"T,
��$i���n� �<ݖ;uP�kuYVm��Ȼ H�16Q�X"���g��LY��=p4�pٶ��#�~#$���gX31���� �nH���K΀�*�^T}�z��.%��&��]vl1��3Һ4��#��V4Ɓ5ҫp��1����� {��\� -��������p�y7OKM��5v��H��'�P��-�ݡ;Z�b�F{�N�-p��u:�8�z��e��p��W ��7`#�r��\Zy�'�����+<�������,��0vdADO~���"��2	w�v�?�F�BF����݈H���y��3H���CtrB��\�Q�U"L���˭�l>�!!Wa;�G���AŇ�K�B�4�
��d�7Kf:���Ň��x����!��2z��fw젲^ɔ(�3����=N{߭?�pK֥E�����z�k�}�����7��`�|y-�~�"^j�lBIr��\:'%���J�[z��ȭ�3�|( v�@I�̘�L7����P2��VQ:҅�@�X�V�
��u�=d��d�a��j�"ڔ~�<��ď�6�5NzV�� ]֦	��]m,���»�9���o�4v7/��y�5T��z�M�xԵM���2��ba�� �v��c��ٗ`A���_ H5��{}�X���|���x�3�yV;l��rM�����:��(�ı���>N9�I��l(H�'��3.�0���V�L��
����}(0��81�&�)&�R�$��B4N���P�@z4V˦�g�D��ڋ�<�{V���S�u?<���
gV�3P�YN��0ּ6�L�X&���@����4�Y������!����%�6e�)�-�8����IƎ�[k�D��yQ�� Xv�Q�-�<�_gaF�D�v�:��7|X������W�Fv&%9vA������2�����Q��ڵ��=ѺI�LmC����4��9�{�u7��8�@AX��ۻz �h�Z4-�ᔨ!���$���Ќ�
[�,t~���EF�M(�ߥY�rH"o�f\�~�V_���?n���; ���rO�7 �o�6~FU����"]��4�S���	�=���,U��M�WVyl:��O#��v����f�GM��,�X��y��>c�f�0�l���XI�5���Ph�%�2 �1���b��R-=��̳�_�*�b����
��h\��[*��FjV��L�@(Ʉ5"w��A-"�y)�{B�HWR�r$ϣ@�vF�|�?u�KI�ӮY��$��!p5l�d���3޺��l��v�8�wx:O����E1��N|��P�K�����.߈��q�N�޶���r�o��b����<�׌�f��1�{�����pc��I:�K �DYu@Du`�B�/��#у�D}�`���N�b�Ϗn5j��G6�~�3�͊o�at��/m�B���_��&���+��6z�~OŁ8�(��o9����S�R�<K��}{�㩓��z2,͢�R��.�z�]��ʋY�s�7�fX�a�j��fx5I�lx=�L���V
j#)g4�Z$��h˶(ѻYF��4��mƨ�Gأ��
b��`���\ו"P�+�����09$Q�c����
(��`�ε��fA�}��e2M Nɘ����?!
���ͫ��WpH�O^{ա�_j	��Od�C ��.T��M �ն��W����G�}E�A�2͊�� D�7(^��Y0�1q��f����!]�_?C�Wa�b�����y������7"ōl<*E�e�\�gR_؅�F��nFL@�f��_�ۦ�4�3�'�h�8����w�K�n�g������uI�R�j�֣�X���0[��V+E	jn˅�oEB"N �捦|Օ�ki=�l֖ct}�� �AO���*�ٲ�� 1U�h�FQ1��l�H<uuAO��i�}���&�FH�V�JrMǸ��x�@�cϪ�K�>h��%.�Q�.A'`�kZ���RQ��m�\�l�_R�d��<:��+]f����65"�l�k�XR8.t��zɁ(���IZW�xB�� ���������_B���C�Ņ�[���~4�5�1~�\ȕI�2��K�0�#��ڸl*��l"P꿤�`�� �7��A���Ҹ�NdK� ��MA����g��k�RkV9׸i/����[l9+1Ff���.'8Z.��ꔡ:[�@�Q����>��C�� �	KVM���Y4P\����߉G֡Rn��u�?j}Zܘ�uF���3���)f����֫��y�j�S�L�NޮW�u�ka[� #��6���S����ƃ|(��=�k������nZZI!>i� 0�i��� >/�̊!���K�z�-����!�_Q§�(��7��r�.w�����}q�^$Vc��Z��K!�?��So*�}XSH�������#n?�H���f%:���:i~�3>b�3�y�v�bD���MD_ϟ���nD������4Y���~���4-4��KO�-����c�+�P~w��tۥ�n�=Ǐ��Xp1��ۤ=^6"��|8�#���Ɗ������#'ʫD=m�u�Q M���U��rW��:@J��A��Ih=�UD͢tM�hMC>%՟�8�c�+��y����Q��A��) �b��K�� m1�1\q�vhX�7����gW�N �!�HO�zv�e��=������J7,'��&��n��hF0i�g������B�d#<��X���d�8 !�)~�a2�k��w)�,�ƃ�31e
�\L�>�K��1T�/�Tq��K
`�֥��B�e6�+ٱ������'a�B�-IGx��C9d�Z�j��!���˓������ֲ��G�g�b�PB{��u�~��y�� �Z�q�1�)gH��kfA�S������?���l�����jq�J@�￥����&O �`�pF�z�j���z �\��j/NB�q���u�����Y�t�����^�h�����M�L�m�2��H��HN!-��k'O',�P����0�-���I֬��RS���]�x���?n,E:� �sy�2�v[O�Cg�A��:
�3������i��8���&1l�,����3�����u���	LU�cM�AL�+qKkj΋�3�I���.�&��r h{����4\.�ZJϧ�ė�αg�i�RP���(<�����x�G��J�:�����=�u�@O���`��e���w��F���{BK^&�@*�ĳgS���u���'U��b�K@X<��@ѶU0��F5���p��ZQv
l���g%��ڱ�"=��J���Qi��7ݰ��:afE�����pc��.Kb���6;�xQ�T��b_���r��)	"��>��hO��Q��#�4z�3���w���scO�.�iͬl�f~��m`1��:�?�_f���fso�t6�E��n��B��L�V���u\�vF�47���Є��?%S�	?8܉z����T�����q���@�U�Eth��x4�g�lM�{���h|*��x�V��ScM��<������d����C��/�S%}��`F���ԅ+}2$���3֢�)~P� @��|�x�>�}��]��_t�� f�=Z�����Hɜ@�F�p@W�%��%��&�p�q��P��d�	ͽ�yO��Ư{D؄cG<���o�R�ty�>/H��|أ]�RG)�Z�cu��g��u�y�c_q��Q"��!QLL�	
L�����vX]�%~�����D�}�p���B�M�:���& ���4�˘@.h5��Ǹ��P����i���W���.�K���ZN�`e;��(�0�tJ. +�&|�BV�2���������<�U��[���l~�ӻ�x)�	+PQˬ�y���W@�?��3 �(jb��Db��Ξ�;�P��'fSG|��ox��53�fs$��G������)��@!�b��d�q��U	c�%��o>]��N2�ZUF�d��M/����X�L���� ���}c�3���O���5�F��x$�a�zC���:����h�\�b������?���(FZ��6��e7e�}����m8mi�.Vf��f�'!G�8�X���K��)�!� K�T�'[�v�%] ���IJ�����6�����a*bRVdi���~
��ײ�ZM�q~�Ta��_,��p�سD�(��ȷ$R���������[�~�7��G�(���7a��ǋ��M�Y7�Ф�ʶ*%}V��T:��~'w�*YU�0����p��W+b�?�v�(���0|q�iK��1;��,�)�E�s�C�ҍ��&�w�q���sbĔ���zſ�BdGV��E
G�J��G�W���I/0�H~*���)�o�=n�h	w���[cTU/�YG����u���)�<��HdAЈԭw�O8�G�P��#
�����c���J���b��{P,Xor\��N���x@�3�Y���د�h�'��f�ΰ��.�hZ5��)QtM`z�E�����Y配M��6@lz�Z��n��7'����d�)@��в�Ls2ݐ΄#%o�o/��\C�Ԧ䔮k�û�t��6�1"��@�k�q�)��,*��q*�h�QG��.�*�G�e�z
,��W�h"��m4��z��/'�{�	T��:$ѳa��2��2�wr%h��N�L��Vg���b�X�hb�A!W�p� �7>_�<H�K@�X�Y6eX,�z�
�*7�ks�t�b-8v�}��F��O�8�C�I�ǜ �Ȣ㫂ۈ �8ii p���E��?gg�[Z+�ބi�CfA�c	)���9l8f�K�D��i�Y�C�9FI��N:�/s6����K��L) �
;y9��C�k��I/vrc���5=u���w�ʥRχU�[��ə'�L����t�t�('�-�>::�M��1`,��CH�
����Bڦ���Z��K�-Ĉ3֮�)�N'�쇱Ă<k� ���#����J�����eHC:�Y����Z|�H�W����T�U|̟��uw�V�w1A�e@9�-=)5�������#�j�W�s~���K�l��ܩ�&�
]�B�z����;Ќ���x'�� ��=#p~�C��]�b��.�+a��謽��=�0����q	�A�a��[C]���
YsvRX&1���Q	t��OǴ�vl��#��S�&K$:Ju_��]L��8���I�aQ���!�U� ��hT�b��f�][�C�p�������Ώȿ�G�%����*��ͬ�ӘϿJ�m�t�̣(Xj ���E���(���ħ�5_a]֎nJ�dp�(¿6.0Z�����_�y�w��v��d��+Z�Y��m��N���MP�o���A#��߆ �u���a�ء�����o�!b���ŏ��� <�.1�)���.�c������S���Z�zui�J��Q����=*�Z_��[p5��ǂ����h�h̲�!זl@��'-yS�������Q8�;�A)|^�T�fBV:&�I7Wo���0vǣã�Ƶrm�1��N.bp�Y�.�x j����=�T����P	4��#�Cl%�F!� ����W&m�U@셗���B(����,%!�zN&7�߀K��º=2��vx��f��81V����7h��KbΕ3��x0�޴0��@O�3 �qʡkܰ���%���\�1�=ʽ�e ��.'���ǒ�|��V�4����z��Ʃ5�7,�2�'y~-��:�곆������8d�ꇯ=d��U�[�@e�'�.P>�ҧ���T0���~CE��=.'���X�j*���R�Q���=�w&��D�c�ú�3���� �j#0�����(�<x;�[�iұ�"��~�BKr7������Fn�}�f�����b~��3
o����5����amND����X��S�[C&��wz���C�.�c��[�npɱZ_�qV�R{��j6a�M���(�iSA�<�؞=�:�)�[�M>!PA���c-q�����J�^pR\�C�;���գ)��nw$I����ڣё[װ�(�#H),�dC��>���&�z]���\@�B�<'<k��<��6�5�)�Æ�;�P�`-�{�+�c-�ny��NsԵZi˅��xlW;Ae���k�z��_C����m��3��g��#�V���
��_=L��nR��(�[y8/����jّS^T�*���G�"� �B ��/�#!�
�#߫_��r��R*V��2�m
�|h{��5�y�qu�k(	�f;�c�J1���\�T��->nWW� ������Ǻb`��`]�@�N�-I��%��	P�w,c����]^��n�*!<�jEa��`��<@h���`��F�������ָ/B�Y�M2�f�Gh��]�f�d�%��Z���]2\�� �>�#�j�@���=���!e��Q=U"��j`��,��+Z�H���`ש����\����,f�L'���㠸I��y-h��P{)n��@�Ց1�:c�79M�����FnB7,J��\���sQ:� ���ⓗ.����E�
�F^ѫMh��T���	T�q�^K�v3id�.�#���,B$����[.��0�����ma�I\��j�`�03Ф 5���kh��������H}��We��T�2���oR�j"&�\�C)� 3�ۼ�x�땪aF1)�,�>אO��8��C�ۊ��#u�H�|j���$����=j�I�#dJ`�\�w�>�Dļ��(b)��z6��L�3G2�h�/{H�5�)���4���eP]-`H~j��X�`}AH
ӗU	��@�^E���ߵ@�A���?:���^�$�F��F�ӡ�����O-SB4jȸ�/�&����X�8�g:�B�fU���@����M��usd)�Rz�{�hMK-�4��J?�R����1i1�qή���E|jS�����+{uj���X�"U ���Я:D�	B��vc2%���g<yRF7_Y�b[h�~'��� ��P����ah	���Wɹ�ܕ�V0cbđQ��$|��!�{�_�1U!+Gu�X��z5��W4۔�̪ĮZB�==���A�#��ԝ����2Pp��4���y[�[��l�I�Đ�ʏ��@ya���8vZ�Y�Ua�먃eLQ	rW����`c��$�@��VG-/4�OZ1�΢IGV�Z�k�0��t;e,�)�1(�+�u��N�?�:ЌW/��A:�u2㧌�z~����9�J�� �C�N��~_x��� $��B���4è��OM�W��hP�_Y#�'h�o�Ϗ��!v���K�<��׈��@փ���KU�Y��Ò�9�A��\^�)�k5�ǐ�ŵ���Iz���jVF��
�eg�@�9�|wd\z�?�,�b���a���W�§垘niu�����#u���c�9���� jc��������x��� گ♗1d��oƥ�N��?�J��f%J}�P.	�|�L�B0�lh���0�Q4a:EQ���$�Ȏ�6���	����Z��|B�^`d�L�������4 Z���.�č�s
��y4��l����4+Hr��o�>�rp�K��	�Ե�a���T��VxC�X&-������CD�a�y�ϥ���*3�On7G�!��J�|e_��]���?B��3:�K�:@��wb�Ps����c13�-��>�e{fpS��C�6�n쩟FUH��b1ꖪ�>�@7`x�e��E1�:8<��Ƀ��$JB�>f�#�֮����C�2��a�*\w3-B�J���g��F�R, �$:՝*�Lot,3i,��2t1��3���PL�$�	�O�㢢:r���������J�iF�	��y,�ML:�G�=�����t4$��D]c-�6ԼnL�r�F�������n���j�&��~�%{T� s�%�TUemWD�@ɣ�JM�H
��L:�	�uO�z̅��Z���@��T��X�>$5�Z�I`��@EVZ)��"`���<�r7���M����bR;�4�Z�To��q����ǈ'y"��L�Ǯȋ�ۀv���2\+%�8Yh�t8����y�:�8�o"��g
3�nPw��!&d.�09�]_X�.5��������`wbt�v�UϘ�����[��M�S͂�
(9�xs�l_$z~��SE�+�-� p�퐣�L ��T9�t��8�WŇ��H��`|��=������7��t������f�'ϊ�f�e#�"�&r�,���7p����|Ǚ�a|�y
,��$D�y���������u�<@lc�E� ���Q�a\�����V�� �Y�J�c�����t��b�u\h ��c � L�Zt��z5��Mr=b���Z���KSY�s5MH�(:'Ev�l�Q��P���C|��55Z�?��6�P_9��	��1XԸ��.Σ�����b��H!u��@1v8�1���~�~Oz%� ��L	8@�x�"�������C�����g4���X�|Ҟ�%��A����o�0L�3�Y��Wg�XOQ����	�	����%�~�~��59t�?Ɇ%��]q[��G����+ 2����_
%�T�p�����lKw=7���CA������z��(�B��x���+�\qb 
6;�%�<��x���q��9Pi4�ʾ��������)ᤡ�b/�lE-��Q$*�E�����B���稿}�q)}���
�"�K��þ]|�����i���V�>6c��9ݑ�H�,e9�@��waQ�M#}�Q�]�����5������?ɺ���෗���I����5FX66?׸����Qh�1�
hX���u��;�}�_Ϣ-��Ə�c��2�;D �����*Z��P̹b�N՜�#�����!�ȐבY���\��Lx�\C�z�A��
�_%�7�,<��
��i�ʮ��gJ��ɕ��n���8-�[���c��k�D��U�C��2S���ˌ6���Fs��**�폲�ۆ}����L��*�GQͪ�(H��30_��Q�����F.�S�������H�<��<9�>�Ϛ�v��۟���ڂ� 󹒲ڞtu2��RE����������c�O�۽����ᾁ��D��te��O��b���ٽ-��i�)*٘����Q�xG�~�q� y��mo?.�o�z��pz� G�i�ڪ��e-��q�y�"��`���n��:G������D#��g�X5M�<��Ͼ��4�L�`��	ʕ��HXwG5*�H����FQ_i��F��<!�
Ֆ]5k����S�"��M�4�rD�|ϻ*I��ů|�uy:e��{t7����O�󵜏fZ�T�8
x?vf�J$vK��T��S�L��۲�4��|�����S͐`�+A N�;j�-����ܓ���k�z�^�P�4&�r��ק���-#$,�W5(�=��ށp��l�]�L㛐�/V�5��{����|zx�b@*||g�t�X3��~�x�p���0���.;v֔M3��1��Eb}���zz�Z������{2�:	�:+��1����}Z^8�Kŏ��G�n�Ż(͢��{;�r���u(�.��z�V7���6�3�Ӑ(^��А��R��+W��T���'���3n�!��i8'S�������	6
��j!�q?9ԗ��d�[���K��K��-n��	~��Ǿ>��&-�jd-��a��H�kN�6t�_s6@�I��<�	�0D����1���Q{t���PT�WA��z��	o/�@�(����f�c^ױk�����<4����a[�/��Y+c7h#6�t��:/O\WP$}�݌�7���oRb��+D�n+����k�b�5�������ݡ���D� X���b�j󇢷���x�m�H!ՙ��O� ��I����s��e
5O���׽��$?��Z��>�S�^���H����pݢ��8ImM�"U�.��3�t�C��S���C3�bF��[�N�F�rǶeD�@]Kq�\u��@�d�i����#�+S��K]H����)�����|1b��'�MfΫ�=xL)�S�CXE�	
|�A�ؿ�`q��b�5F*�C�v�Ð��
W��|���-w�q����#�؞�ɀ=�!�
k,��q]Oc�j��1�ٮh��j�U=�}+F��p�T5��ȵ#��s��;�Z`�6�x���uf�ն��OD�"�䋋���r�@��!w���p 2
�w<�O�Iw9=켷wY,|6�o����uol���vsl#��L`���C5zʑ������⛧O1��J��D%�c�N]��2�{���7Q��8�"��PI�������Ҁw���8F�= �7$��p�S���^[�������7 "Hd�o�	���i෉TE������������4��À�sw���~��5�M��|F&	�Нh�n���~h�x<��3H���=���X�(@�Es1�v ��^?�����(Q�#����gՌ)��s�ؗn������#���m܆��ouTݠ�o&�f�3�(��!�h"��ȩc�ڗ3��XP3�͓�i��H:��J ����X��D�\6)�(j����ıh0�
B�W:�]�+~n�8�k���2�;CM·����{�ÛX^=����]�pzQ"��xlP���`a�2@�P�>�t��� /űx݆g9mx����#Dm{$�A|NQ?�t�ؑ��l��\�W���?⒴s�XtB{� �
6�[p���p2�p��ۃ*q�E�e�*�e��w�N׀�<��Z�>���I�ht+r�����������u��|�yv�8B�0}Z�^�Q�8�a�<�W��y������_H�Q����qЋ��X-�ە���S㔞,��.�o&|.gKrP�!4�؜SD�Y9���p�H��Ml�"�V�E�f��!�,�٢������ZƜ8��4:�x��#��VX]%�R\�˫�� ��8�p�3��)]�#*T�&���㺀���t.����1�|�b��4$�8V�L�؃,�KJ���.z�ƅ�Zx�oӖT�Q���&���y�� �30���9W�G��*e�:If��fa#ۺU���iKVɲ�]�_&PY]��97K�l�`걣o�&f1���ٱ����A�f�`�כ���BP��n�X����7b)�u��P�DD=�n=b!�vG�m���5��;���\��g���6�y$�Z���&���@m���0����rP��O
[5��8W�s���~5+Z�?$/SAA��=��t9-�s��3�x�'��bɷt����G�<�]�LS������:�*��� ��:�b|C6����c�2�de)����Ӷ��@H�6;C��œ�' �p���|�{���DTت�_�̫�,ٳ"N/���c,w���b��Q�پ cB�B@�3��7�i��� �C�1�p/���O�D�Ĕ��XԀ`p2T%���ZƊXǥi]��x=?H)����V��~[�P�d�C�E�ܘ�%f� �R��1bm*V9���b�~���5,��[�������g_��/m�n����3����U�]N��x�&d�c���2�Z%uS~j�3ޑ�	
��pX(uq0F�E�FJ"H�O�v�!���X�_-gd��f.�B���8A������օǨ�C�@���ǟj�_��w��Ӷ9�SP���u@�,�j�)߰m�F�:�ԀV�!l܈6��� A.Y��ƢԚ��ԚtN��
����� �l�52�Ɏ邚�蓗Ü(���g�=�v���d��p	T����u>�ir='=ԟh�hP�j�l�hFbfԭ��~�~����j#l�Cnq�ή;bͻÛW�B��t�������o�E��Ȓ
!&�0X^���PW���CA�\�4�iu�M�8�3�,���ϣk�J�	Wh��K Zc��;��b@(��f��Wb�+]Z�0rDmÂ �7bw�h�m�[��	������_{�Q�&��1� Hb�* �� _(����I{���<��1����+��ے�#"�RF�z�XX�&:�w䱌fGkVW�g�3�c��HϏ����U�Lz�_�C�ʦ�ƞ8F����=D�e/�w��[e��0�:�$��Л�C��Yh,j?�M|)n��>'���Kf��SsJO"H ���C�)C��a��oj���Ǩk��/v�q������r|��C>�;��!f1?��Q�)��������c/����e��W}�u,�s���p�㭺�#�k	桰���Z؏c2�{��)L��N,8���e=b�F%��Ry��b���`լ�X�p�*��qo�)��پD��ؿ�H�!,Fd%��7������u3A*>�o~�`�ly�0�+b.���xhPZ����aٶ�W�oA�q����D͓
�T�/zu���/_�����Ò�y���*��e��qJ��j|�o�
qF _Κ�]U14����5���=򜰱� kO�T:J[Do{�h^,}4Qy������{f�k�sU�&we���`q�c�LH����I�<�j������%� �3p�P�$��=J��<]�/�[V-\k=��p6zoU��?o�A	fל��u�����A��/�
��i"����/ԩ�V�G�R����8UT�'����y���G�F���M�