��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su˸Y��'��d�Ay~�`�i���o3 1&����1\T�����	��!mF��
��\�ݘ�#X4|'�~a	N�1�""rϗ��?���ݝ��^��lt����d�k>O@�0�#/���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>Q�y�`�}@#�����ڽ�?��^��'�eO�K}�:96���/�F����+�BZ��1�i�I���WLuY�Ɵ���
�g�(q���������	�����ҁ����)'2hpf�t|��нX
#c��7@o$��Ȗ�����z�5nЛ����G� ]��ד-'@|ٰ_4'i㻕�=D��ϝ�W=��s��aa����:Dbޭ��.�����m�Xd#�t��!��4�,�C�����QD��/���1P�l��/b=R��)E���ٱ�H���Y�0$�x��2�*���W~C�T4V�pбŜ�����rTD�q�Y��J�(�  ^3����h�1Ս�٠,��ɼ�R�t��H�U��e=�]U�uB��\d\ϳu�>��͍�~���i�eE�Ԝ�#"�[h�WA/��ٶ�E��N�Q�=����;3���=I���s�'�A�Q����6`#f[��کr��}_G��9�Mɶ(��*�di�u*B	N����"
\�>7�H�q�����.��Կ|�J�x�q�X���ZG(!���������=о�5�d�DY�ǩ��|q�{4M��t"@h{��Y�p~=�����Q9���F� ~�-�0��,��^���۠�j�E{�Dw	�g��x�ȳ�Q���pLx���s������%�
�s�Y�M�8�Ŝ0u���p�QG���O� �.�:4��բ'��Gr�=X�` �7/��nU�H�ɂ�U4��ƛJ��/�Fc�<$9�L�<y�Yh?�щ?R����6�(��>��q�U����$�U����J��7�lW�JZB�җa;��cIh��^"��q_l�m�ΦI>�����Y\��MmO��/�`}q�z}a�H��î6q�z�ҟ�9�vs��L+:�)>8�m�9�ҭ��� V'=�TK�"J���oB�K0ō;����G&��;�������?��&�ڀ�3���4�?�.�|g�E�P����N�9BS��x�6?�N�x]ŕ;����-J�j��9J��^+�C�i�*������Y��J2K~z�p���E��~>�4�)���C�κIY}
�^kJNN�|�Vd��d1�a�{K��Lh���%n����x�~��_��8�����u�,�)�RK_/�oqOõh�2Kt8���Kg��U����rF��'9��i�r�o�\7��n���)q$v[�,����:��"$��!g�z6�˙���7���ƓQ�W�`�/%ꎦ}�hՋ��5�/�i�^e���>|ߖ���D�3�-&/�F��`O3>a�8U��,������<�-�ޒ�wyy=�g+I"��Ws�N~�,��`4q�8S=@o���8՝-5NԦ���?d�K�g}�I�MU��a���>����3�$��@�tBK>�\�B
��W�N��|;T�{ ��|f�'�E�`����3@먂�%������`��y%4�Լg����*7���oʌ<b�j�*1�%�* z�%�hR;5G�	;X�!��Q���A�x�jz%>$H�r���Q؆�L9�O��Fq�>S��F?��w�R�F׼����v�Hdt m����^	k@�tY�&Љ���!3���Ȗ�I���CIt�`l�M7������4F�(���:#xB:�ǋX�-a@�\A҅��%�"������M�P��OC��`��|�|S4"��B6T�� �������&Gz>W�Y���^u���r�ƍM3?�lA6�^����C(
h�v�յC:����:�7	*O/z�d�oL�]t]2�I�'����@7�ѩ|�:�fь3�d;�k�Dx�&�h�`+�mH��-�#gAN*"	'��9�U���e���e �*ء�1�5L����ڐr䀦��/,K�*�{�>�t��E��棚��'�*c��	ۗ]A����xg�I�*M�$<�ޟ(�mb}�~ЦR�\�c�K/�^�����j�WN~|��B�_C�c_����3ƕ�+�K��=��^�����{@�s0Q�Z̜׏P��33��-�2r�%D{	��A5��u`�������F���q1F�����Nydd�v-a���S�f"�Q�~��P�@԰rE"o�����J�pJ��1%����U���k�L�L,f:NNNx���lu]ؠ��x�66��,h���2)��U����d�
D���غM/oi�~a�@U5�O/��P_,'/4Y	t[UT(4DR��o/fٟw�g��������'{��J��+Rx�2��u#�Gek��\|������2��/*ㄠ�:�D��%�
P�;�K��[ζ�*����^��/���K�=-���Kl���L���9IS�St�'ɛM2 ��u@���Fªb#�9�Q�����X�ܒώ`9�QW�8jm��&u^ю 0��
E���­��o�u�Nދ�ԶȓR��ԉ���b�����fV������t��H��0�م9a��\k6qD�#t�K|=�=��a�X]0�UTG�We(\�CR���F9�y��blkb�$�^���M���-]���Z?D��.�Xo�A�+N�9A���������^IY��+�:L�Ϲ��'�ڠ�'I�ptt�3��^y<�ǈ���p����އ\ H�hʘ\�S���R`�|��&���%a����D����!�W-��Ŋ�GE�ZL��6W6EIDR��6��)#��&0�/z�w;��҄���>I�5��Dks(K�T����|�9;'k(��s	ݘz/�w���{I��9�g ߣ�tp8�և�Z$�Ǆz) ��)�L�X�vU8&9(O�� ��'"���@���U=�d��G8��]���K���l�Ͳŕ
�]���0<^�,���o_��v3\BS�>�څ��)+њg<*��n�g��bL�Z_k��J ���qڵP̀������r��Ec���ZRr��0��'׸��������o�*"�)o\Px�� 9;�$֯�EP��L�}�+1ST
|��'���卥j���X/O�qL�,ʤ�X�<q8x�<��R���j�+G	�k�֚JL9"`��8-Zpe|#���ޓQ��FT�!VJ{��]akrt��15���;�3;:�/�c18����4(�nx�`}���Q��'�cw�햗XNr:��u������C����7�̂����HoI��z��{��áEfuf������6��CH��;쌳5��������&��A��:�t��3M�Wc'�j����BH�	���SLR�T�]=쐢�9�D���3í�+��1n C=t���Z<T�W�ej��N �v�S�ړ4W�Rk��u���sB�+`����0d���ӎ����/e��I�����ѡ��:d��I���	��i��T����������h�ݧ���zUB؈Fa��0�1^�IuO����\gKjBrIO%_��ٲ-��Vu�^�/�Bو�y�0k/sJ�|U����mm�\���>�f?��	T�Y���g��,���K3�%��^˕.rb<�j��5��nh������V����F`��o�a#ڤ@e6�/m� ��FS������t�֎�􈛺,��S1��c<u�{����Ώ�ѣ��Y*{�;�PW���{	�=�!�(7 ���-�	�}�%3�@YUȮ��G�i��fT�9�\�J�R}�<��!�+ę���Y�/uخ�>�x�5�5��2�@�6.Zv�{�2��*1AibG�_���3K~wX�J���`�[8Eq*��&{�"J���x'įE3q�s�}��ٹ���Zւ�|�����EX��/� ڨ�xXҸ^�u�Z�K��z�i}�s���K&<W�kA]3B��4�n�<���j����"̥�@l�n�g�/h��䕮NN�)8E�\A���%�������%K	{y_��
��t�\�Qk|�ߟ�2���L_C�׼՞��6�`*�Q�Y��֨:.:�AD�d�`��ٮ���`]��W�<<�c�ǘ|���D3�|�͍T�z\�|s߱�D�
��y�������������=j���.��GN��v@�y�*Bb�`aĻ�t^�0�% i�����i��F�;�׳��e��l�����#��/e��>���mc���B�� �l��<�2��3fC��1CBH��2�%���^>׀ؽ�%�0�;�,��� ���d} �����:���sH���}*���{_e��IO�+&FH���4�g�<T|-=!�D���C�:Tb�'�a��r�2.�HM�20� �ik<���Q���R�g�������X���㱔���>Q�E���h��0���F1��o���-ہq�`sR�g�ڙ��Ku?�z����ǥ�~�6/��Ku� ���4N�ǿ�O�pv@�q����5v0�F�QA��[�0%��,��N�P�gV�^��������n������A�3����mV��E��+�k�Oz����r>�InPz� I:�Hz.
���RЁ�q?����\��a��I N�F!@�� *k�k�E#nd��'��E7]���{��Ԣ�4B1C�)����b���Uh�A�X��>�-��k�CfTY�ȉנ����dy �!r�\n�ٺ��!Sdgl��ʰeh�a�۫8Qޝ1����0?�;��KH_�N�f���Iu�A�*�?��/}�^
Ϻ�"aҸ�_%�����S�	Ɋފ���js܈��C�%���'�[����-��J��JhJ���.١�t+�/��pEA��9^J��`$���/LWV�ݼ�0����k�J\��:M]QTϲ
���7q�F0��k�&���*w�5s��{Yw��0�t� �k�x���Gb�g�45�	$��Kҫځ������O�>��g��X�XB��9�����Kݠ�&��7���}�NZ �.x�o��t�΃*�W]�D{L�����Z���&i�OH��F% #��f���W��5p����y�� v�%�V��-W8��ghj׸�7�).nrAlE��QYQa�HG�Tr!(O��C��µS��������O�g��=��H@1�A�vІV�{�G���t��J.2��*S�88�FFv�@�����-����׳z$�P�����53�`��"y��Zr�ɉv����R��n�fͦiw�� ;hڥ�yv��;�M�.ԟ�K����;68���]�Z}778 Y����7T3�äV��o�E�Ye������;tIJO��5
�(�7��v����`ꑍ�~Nr,p�.n�M`�h�1o}��HA�c}QN��;H�q�ML�0�Qu�� ~����	XRH���`=>�M�H��p��ݨ �`y%�Z�6QȒ�3���6(�t��Y�@��\?�������͠Sh\�@�Fvj�f���'k4�{.�Sm�zX��p`�I�{���gs���T;^�*�?�*Q���H���q=��ø����=�DvчF��΅dqL���3�Vh���hY�K���i�٩慕�(�2�}8������a,��Q����J��V��(�=3׹�Zj�}R��b\=� Ӎ�g�4x���M�4h3lظ�((x-��6X�9;�
4�U�
�ӴQ%/�&��Fj���ҭ?�Iׄ��f�ɿ�����,�θ�8�ͽ�pJî`p�w�7��T�X��@w�O}N�j��ul�S�e�}��0oe���w�7�&H�3
��>��;] {λ�K��M�;kP�d,�S��[&��q�OsV�2���.�$?��D��ث���~i&x��4�H(>n�n�dY��?l_S{��U��5Y��g�F�k�`b2~p;j��ܧ��hFi�A�u�ɢ�����fr��z�L��n��0~,�uś5�\�y"���ԔJ#��G]���;��P2���#��QΏ������2<�p��1`(��
���_��{���/�F	����Z����;�
�y#����}RD��U�2h!|r�c���S����W��_ ������-� Ly1�Q���$��'��\P��i��Ҽ�-�%*�D/+��Kݏ���g����6�+��/q���ӓ���C�&g��|��&+�w�+|���T����x�X���]�k�%9�c�����d�q=1w���
M��D��)�	�pS`P��|�����~��&;���*=�dj\�������U��H\�ጘ��E]��x��w�1�;!��̺oĴ���I{�?82�~�Y>�*R���#�aV��ӯЈ�)��^�\�k&��O��hƄR�N|;�r 6L�z�LB2\�AJ}���'=�'E8��	0���p�ڲ��2ѐ���$�c� �x$N+-�E-u2�8��L�Ze,��u+7$� ������Z��"1.��}�W���4&	:EL���~x�uٟx�jѩ�5��"oT�3�D��P6�W>�;�n���!���Z���W���C�"経J�l��O]<�p�)��p�v"b��D����I��'#���=}ׄ���!y�|녻����`�)�����^�������_�e��{�0�=��~,�ջ!��}@��F�ǁ�L����:��,��J+~�4nF��Q�{ӆ�;| g6?��B��2�8�zV�IJ���\�ߜ�R#p�K3�.GG���Y�|���Y��+`IO�P�&.DTU���2���`5q6J�VX��fڏ�h���oe�>������]%v�vK߉�ȥ�z��ű�M!���6/�L��$B���վ /���\i��pPTQ�Q�w�_ ����9��O�y�Q��Q���ݘr�j�"c-��T�'H�����庽��F#G�?7�r��N�I>�\>[���f[�1�->��o�z��,С'���pk�����I���ƅ�#�+M%Z�}|��S*rq��S/��ߌ��pʴ� �E*��ږ0X�L�:���8X��P�������dɟ�Q�Sͽ6U���U�T4�39J֓/l�Nk�l��c�뜚�YP���6�W�n�C+h�� X�O�1(̏D��̴9�rH�|�=�ȥЋ�}q;T��SHv�o��Ǌ1��S��B��LE.���D�L���Wo��üJ�k����x��(\�Hf�c�W��?���r���M��a?�	��~�2N|��r��~�=[�>`
M햎�g�'V�������],���<��Ci�cS��	
j�0+q�@m�hǉ����N���fh/^�
*R�I}j�itx�R����S>��oN��</�=��Z1��e����V�4����~�m��k��8�X���<��l���Ƒ���,E���t�oʄ����uڵ�O��������f��8��&�*���*�Oj�ΉqHeHZ)hwA�+�6�<M'W���͜`��'|�,cE ���E��Oi.GI�1�^R�ΨH�|���5�]������=|�ݲg|���y�] F�Ԡo����FF�]��U޾�Q�k��
N���	eĳz/5�#D�x\�'f.�AC�=�,&%hzY��tl|Ц�.O��,�������P��t����c�j�w�r��^�Y��a����+w~�:�7�7��I4��P(��H5���u��BP�a�5�Z�Y`�cJ�6FF�b��N���D����;m����-��x.��^���&y_+�7��E���3�Om&��(7��s�!L-����f��F-;&�Y;�6q	u��ʅ���,���}� ���w���.�܁޵*է]E4���rk���ŎDz�4o�Ƚ����V~�)�:o�s����P���݀��~x�)W�Y�~�:!��d�Q�=>^�&#j�Eo���AUM������-�2y �ߠ���$�
�$Jz���������g���"�q�d�q���.x��8�Ni�xV񒱈��#���>�B8���{�kYl���Xwk[L�%��X��x�ap����m��R`�'d���<#��b���T	}�����G�Д��3��.�����/�(�]Yo'|������H�#�Ϋ~�6�V�Y�7�t���B�2��j���=i��W��2����N�xO�\0{{��S��^X����&}�$��=g�&g��]|��C/�80�P[�&b�A�k�F��{�dy%xo�A�;8y��\N��:k�u�r"7X]U�^�?�Z�����[�O���t��=����b��U���}",i��
����$�2��6���ny�O��2n��&��>��,���h���t��׵�r��`aE����h7�����Q��d'�t�
�w/��Ǣ��:^ʇ�kgv%/��7���ó�[&�$���윿ɲ"�q���E��
��������Vl��'{Zԁ��d���d�2��5*�8(��0�0T ����y �g;̀���[,���{zzI�h�K�nO��/I䰜y"����!f5�Z��Tcv0�$|�S��?b)[�,�-���縏`�i-�a��GEZ�i�����Ƭ�+#�y^�
UK\0�%���@�@�Z$8��eY���m� A����Г����7Ú�@�A�E�?z��lA��͊�C�(6m@ �@��%���Z��$wT�4;U:�����X��Γ��1>��Z�x��Y/,���Y���V��Y�>�cMjR����f���ME"򁰭�>�M\��3�����n�ȋ�rǷ����-f��'g��N�s'�- j��S>��T��L����x��#+ȣ�݅�_�S_�2i����2���?{u�x8�ڇX���I/	<B�&��f�#U1(�,?q��6��:;���+�_�6HQ�o�؞�Rg�M�Ƈ�|��xr��z��e2���۶������{��0ôJ4*X�i%����6[�y�Z��0���9���?�V��d,}�!��9v	�6�E�h���mx�$ҷ�cB[�'���K��2k��Cax&j�(Q���dz�M*sq���J��VD�tG�JEW�+e\+n0s�xMf8zJ9O�Cw<K�b}I�Ī�2��D&��Qz�U�b�Í����!Z8	�=0�rޘ��@"L@�q��M��,nN@��n��<����*}ش�R��W��| e���Y�ܸ�w��Z�?nr�Qۚ���oT�5ϷP�J����"�O)G6���ʴ���1!��&�g2�L���aHU�����Ic��Uÿ��������òņ>t;O4z���蟂Y���5���v���g17�kA��Dߦ�V�&��yxtS�Ѿ
�I���>�	Y�	X��W�$K�/w�;%�K�5��{W�ܕ�%��?#�2?��v�Y�a�d��>8�Y0�0`?�J��s�����p���������,���/��ll�"�2c����x�/�Y��<�2u�����i���3*�C�,�~�V�x�X�z���X�����p_NC�s�"�7�J-d�*�|��=d>
��<�N.1M�����|����I3"�9A�UI�<!*�����C?�F�� ��t�I�-��MP���L�o)�[i�bk�6��z�^�o`׍�W����9[_������Y]�J�|��H!��ق��i��b�P���?91٪�ߝG_�F%܋��Gթ@r,��gę�7Rf���M�P�M��x����.�X��R�H�
�k1���I鍤��Ʃ�_4pͥ�x?%fyzJ����T^����_KY�$�%$�%��/�N$F��&r�P��O��S��j�f�9|�w�?3��.Ԏ����+X�_=���])v�tL�`OG2mZ��*�ixwζN̶|^�: 9d
��޼92�\�ʡ�\��kl���P��cƣ��(���}���*8���pMdʃa],����0��5��cx$-gH/K�R8�$��1{��X�VF��'�E����M˦"�h���!�癃.1O.O{��F�,�w�y�}�MP6��U���[Ԩa�lE���TH����`31`�����/h����5ś��FS����˄�d�y���P�%�]߾O��#4�w=Eѵ	?�\9v���:���uU�K-D�fCM�ٺM`�
��6���dVT�6�gJ������Eu�>�f!U��r���Ju�^��Z^���x�|���S�뫄�ݱO8���P[��T6�[���r�Q�}���dl���C>b*��	*� `���(�r;���U�.˔(l��}F!�H�?�.w0� m4�LNHUF�D�Z��"�g����ʚ�����#��r�3��9{��%e_�Swp�؋D��������{'���id
��J�PlLi������DA�hV�"�u0h�̔Z֤<Wm�YW�UW���{*/�L�w�>�J���lobD+�`�J��b��߻C��tY�!E���p;a������
�����T���q��܋G����v���)�%!�W�8>��"�!?�YU<A[
�XD��-D�1\3�-X� E0+9�9��PL]���Wb[���Xjsu���~^J:�vz����>�����A��rሉadQ�{���}s�ƌ�ct���A|m,>W�C1Tu�9Yłi�0K�4�x�*��"��Y�?����1\��/gRB�NQ�}��x��|ZS�n��q��]�t�|�M�u���5����?^>�.ۂ�i����R�$�~�%���o�kA�㙏dr�9@,�+�#ʶ�l���?oj�j��L����?�d�,�'������ι�^�yT��o��-5��с���W�-�Iy�ZW1����`}�F9_��������#�[D������0=�qV��Յ��IR�d�B����v�͐�H��ht=��B�ؾI��IR=+AE@G;���܅�L�~E���?�7����,N\�o�8�ܸm|���(�:�2���Q�qV*�@x�R6��#|�lb$#wq4�kmEI�S�����O��CձL�I�|ҏ�2���5����K%<lܐ]�#�=s/�v	-�=��-Nl0�EN��-�����ܜ���!��F:�q�H9���#�ȭ�����;S��