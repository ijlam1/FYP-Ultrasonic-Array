��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su˸Y��'��d�Ay~�`�i���o3 1&����1\T�����	��!mF��
��\�ݘ�#X4|'�~a	N�1�""rϗ��?���ݝ��^��lt����d�k>O@�0�#/���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�
���B�+98����E�	�ۀ�}&M�8r���XFT!�a��#��\DTy^�@�tW��\��@>Mx�[���l�Y��/�w��O�V�vB���}�_)���t���m1S�撅���Y���N���?߈��� ��ߤ��'�D������YK���NiWig0e�VHc��0] �f[���Vʐ���iTA�C�C��������"U���ŧ�!b��^���'We�Yg/�<ʺ�=��gج��cңɩ�
����U��cAv��3���L�$G��Y�aZ�s6��.���h�*��d��
���f]{}����h�29U�I�Q��"���\g��;8b�!�om�f����uzXx3V�2�v"�-����/���4����#��'*�U��;���y����12��#R�@�@��R�3�&��q#D���/4o<o�(͕f����]+b.R-,��܄g�+{!��,_�h��R�2����nt!��m��rw���p��c��%2�k����V�CfO���v���e5����8�,&�������� �X%U1��!�����C�h�5Q9��+�b���"�n:�PN~1x+ӥ{�S�g�� ��=-��kH���'�1���D�7
X�<�"܃���&����=�֟�gF���#���n�3�a�>��֐uj��P��N�q� ��قȕ��l���Gz_�Ą�xjV��KF�p.�Yq��$�.���B��|Ei��M�!����������UTԿ�>6�X�:v'�̭%�j�;�@F���5�B�%��J'�N�P����t|K����z)��W\[ �q��ހ������%)0^�)�.��^WI`��7p#�U� ��Vo>D����J�Z�{�UJJ/SI��t�,XH�8�	@}�O�)�HQ���WV���� �^���W�`��@�. ��t�<E6�D��p*�����>�H�=V|l�\x�{A���[\�`b��;����qyX���yD���?��]�6�$gHs:e0�0�x+��P��>Hv�6-Z0�f��l��c	9(ݿ��J�YAp��0m��}'a���p�	(���$(��ť�N���8��[���<�C֫K5d����6dv��/��߬Bm6d��0���!ǎ�����旼���LtWZ�Mt=���k�o�����
Q��e����5LJ5|-n$�'����[{�8(U����!i�@��C?���0!V��B
l>��m�q$��^���X�˴Pʞ�o�I�X����X�n상�s�ck���9����K��(Nhu��=�����a��u�P���u�$�s��O�#W�f������eJg�NT�DX���!�͸� vH��(�ܸ��	SA�)+Šuc	)h�ƽ�����7��W�K��Ӛ���WA�W���, 1����J��esu�?;)�/(!��+ƕ(1��Jľ >t��Y�ޭlj�Ո�OeT�a��u>�H�/�!���6�'O��0<�}���k��L��5|�j�b&'-�j�G\�6�|�IQ߮A[�+�Q�EQF�O͠�]���9�6S�N�=���(.� �h}E�J�w��\����|�%�mZ$�Ǭ��n��[M�ӻ
�\���9pW�L��vZc��,,5R<�ѲQ���70g��H��#�
�9@D-���lJ1I����L��4͹v��g�57��
o��9���>���'8���R@Ԏ'A� i�^}�����lK���+�^��"���4	&U���O.P����A
��� )��}K����L��PW�^���+���A4���J�)cĭ �G��DyD���w9	c�N����h��,��X��Oh��j��Y�|�����P`�����N�˛7�����j��8��L"^۶�.�U�� *6`�8��ܺ�g�VV&�f���N}�����V�]�n����ESf�Sg���k�k��(F�4G�Ŧ[!K�ܯ���a�Zj������������2��[���bh'0a2k[�I(Q�e~j�{�8�KS�gF���<�3���;W���I�v��ɻ"���Hv�%2Ϫp�HW����;a��Yی��	F8K�N�h�[��ڦ�z��3]��4���S�xB���x�)��C��/�\"/����t#�]YYg��HwOϲ����]�Y�R��yN� Su��[BSE�N���-�G(��mT�穅�"���C�9�ݫ��h嬭���NK�����$'���$͝ټ�����s��G�f�ˁ��Y,��� ���lR���@�"B���kD/)�8��f���%�h��)tɒR#�U�a�ͺ%Tt����$)%@N�1#\��yI����N��n����V;>(	�̍���v�wug�)��#z����c6�
��	��� ���R�}>$��j?����@�]C��.�����某cN�x�5P]z�����]�r@!`iT-�ӌU� DN?�d67�Զ��^�+9}�4�G,Zx_^
0��s�E��#v�����q@b7�X��P-��V2�J�"��h/G�����j.<C*f���SF���Z�^��h�6�%�d
����T��d��Qf���k��������$-ч~<�H�a�B�a5���FIq�0=tq�)`��>��Wv��$;�雎2U�8T�p���W4 ߩ�I�|w����Q#�G�~%\�͜;D/X�y��鄣r�W'��3��9��Td3w ������d��%!��z���%J��ϣ�)~����I|�:Vg7rc�.���� �[���ׇ{��7�)*N�6�G�8S��n<t�q��(C)�ٞ�j�=zj��0�N:c��B�l�?o}��(@�(se�0ᆳ
�q�Y?���~Ui	͠G�v7��YP��/�e	o[��W�4���WC�CR���<��}�iM�źa�4���3j�Q���I5dyJa��L��?J� H�`0^b�ܟ20T�fPyd�j�HY��/��2Q��������*Rt�/8�Yv$
�8/�W��h	o8�Nj�8��Z��i�HSh�¬�{O�1��4*���W�w��A?�o{���4$�������ă~�H* ,�>F���[2H��>1�'����xR�Y^��n���M:\��հP|��nbG�������S����`��d���fr)��m<�z©����",,i�O�Ҭ��TϠ�+�rI/J�w�D���d�}��@DG�ć>����<<2�8��]R&Ms�[W��"��KO�ж �0gH�w{��iԧ\@����x"9a��`���9R��Ys�2��9�B�J�(/��T��EV|D2�>X&��8������P�*��BI���d#vi���Ɛ����|�_���ge|�R��l��ᡓ��J�s�9c���po��G�!���ip"K�����$�Yy2�����j��cf&ݢx����;%K����uR�MXr����w�y�Zn9:���_�ҟ�u�t?�P����"E�FwmjG��)l�Yl�
R�/|������y�,6!��%��u*Ŋ���R����FcvP��G��AY[�@��(w0,�y=��ʅ["�*T^��� ��U�B1V,��7r��յ{�� �D ٭+:��|.�Ի���{G:��Мg.(��oV��U�}� ;gA��V�+�B�y0��{��H��'�F`�&*JӠ��m�R+���᤬���N��%��wv�b�o�5�::����(�J��|Hu����n,=t2�T!iHWEz���G�i_�^F���[횄1�`T_|Se0ݾ�1����l�?���7�?Gi�G�$F۱2�lyY�"�d,�A�W��#\�3j27)�
�nښ�G;�8C�<	�l;~`a��d3@����6�D֥�)�;%���RS
��3���	E����	�١n�8V���`�0H0	X���WgGz�:��p:pN8��u�`V.�Ad�;y	g�]ΑA�9[�֌��ge �$��#~�뤐��@�cg�{�=��#���?�OA\��ΠV���l(6��36d�i��:h��>i��پ�)28��C�����E �E!�SĨfz������p�<X�'���1�RW~�Bg��2�z)��xt�
���@�,#
*N4�;�N^gx��(�Z4k<>�c���Ȣ�J/{>�cPN�vi ���	������8�2b>o�$'������nNtN?���NJ�bUi��l'�%����G�mu5jϤD�LV!#���>Uk]9{j���	�v��i�����F�u�9<���8�#4\^�pB'̌��~R@y4�dɐ�aⰇM�e�>U		�������$���x����a^���*�zD��J}~8���]'�;�X��_���Q'y˶1�g�L�����]�N�ӏi��Ǉ+�m�=<Rܔ �ƺ�P�咣�mH���n7��edL��K�������Y����;�2XBf��+�Ă}�9�����Ɉ�������C,3 � UV�!Z����1����@0^Ò��r_0������A��tSL8�]L�p�Fū�D����,�QAy��$#�q� nUx�8��ULf5���^vy ���z0#���H�=-t;���~H���?fQ�o��*��I��3���sF�R��WQ����W���WSr�m�t���#��=�6���NJ��[(+f[�3��J���/f��r�+_w(�w�а�8��s8$9��8�4���:aRr�)��A���G��w��S�(��t�T��~�
pf#��L�H�;�Y�u�KÒ�M�۽:8Π��"�ե�B��+ሴ�{��#S�Ut�)+��ę�IƠ�t��O��M�*R�z�[��q�T����I^4T���[�����ap�ȱ4�͉�s���q)��|���?H��9i����r���$l�e��&@�w�\P�zۗ�6�㔶��cE�z@�N����2ɬ�3��#��DF��T��Q'&J6���J>p}���wc!ǿ�.s��e�!��Nҵ����jw��()���92>`a�O��QCȢ%�O{�HQֲ��9��M��D�­B�t�i��Շ8����'EL�p����D8v��GR�L�K�>�%Du��6!4�f�&ˋ������E��w�Yeg)��'9Pi�*s��fh����#�{�F��k
�c?s%=�_����;��%�b�iK�s��q}������{;�f��y�\C:+�t#�M��reC=0
�׎е~a��mޝ�}s	p2��?���Y3�*d�� �=(.��cc��9Bx|��+�#s|45u�.e]�_D�P�&�ƃ������D�Q	��O���R=2�	7{����P�Yަr,�*���рl$2.ˤ�X�
���$��zE�3��2�5s���kz�	��4]/��=��_,{J@_�\�r���LO��:6:C���'d��I��uY�`Eڍ92�L')n����,{���z�*�+-�n��w r_%�f�I��?ړrg.�����LХV���7HC?��P�a����Z��GO"m�*[�#G��?�?�i(��������]��r
�����t�.ذ����}~`�w� ���i��d3�v�%�4J:tZ�Ak�?��МE�U%U7$]��
yA�]�#��"|��Y�d����|8t�~9`�4\@@?T���H�S�(��P�΂�Q����9�ܡW����fA��g�����7��a�'�͌��b�1����t�+����_y˾cۥV)��^����`��4�T0�<��ŗ��G����}����=�M6��:��ː���籷(�aK��~u�dD�|H�n�`���߱���ɢCN�(�>:G/ ��~	T���I�������QS��ǆ v��� ���A�ݠ�NgN�{�X�rǢ��jʀ�p+��E����p���mU$��Վ�a(g	�����_UH�E;��(9���Lb��ӥ��NsC�c�ݲ1a4Uƿ
���������X��d�
v5-b~����k�T�z$�m6�{�rin�6-�fၣ䨖��Ձ���y�^PK���˳���f|9����S^�pM�|�E;ƴf�Ô�b�7��T)����2$�>�6��4�)rj��e|"L*�^�	��[ ˺���LG���9���/ ��aD��;3���rz<�R�X���=��˻��*z�1��i���}���*�ԆexiE]c,4tmO��sM_��bI��mL����I�)LX�*���YY��'(>���a��&>��]���������<���СD,މ��	@�sҐ���BN�')g�J)Ƹ�L�]=_���w2�a4vQ�i�e7f�nM��T�?4�H�u�*8�G�`1�=���l���%�=S��)w9!���S�?A��OȃĎm�Xا�����#e7����|dGq&(5��D>X ݟC�ծ��*	6M����J�)\rC��h4'|�����`VH!���?�?�2�i�|,g(ni�p��:�k~[�W��'�b�����u�"zh�Tji��Sn�T3�pA�;�d��v�Wܖ$-c���+�j�W쐞�H�M';�&q7~����x���.��L;.�D�H�Z�IR�J��_�=qic^˦���=6NN���WO�A:6�B>jKPj
O��3��M��J5�w���J�����i�ө{��Z}��}�&R��x�>|������cv����Z�Ԓ��-0Y�ҝ�+��r�.G23���h,�֣/9Q}����珳�|��.��^�`ܕ�;���FS���}7M�@��[�Od|�;�l.�Oq�	l�� �j�X[M"���kE��R�9�ָ]�V����GBӴ��f'䟏�rJ�g��}u�Z��N2����#,�$�#Ox�	5Ʊ�����\߲�I!WC�aAڜ���=TS���ʦ�~/ѱ�����ȓP�ɏ��9j�<�z@pbb1󎆼��������/�>���=�d�P�ŷ�Zy1s����ͼQ��~�޹-Ԅ��o17�ƭ�0�����z���,9�cY"����I�a�1���<Vn��c�J&l��r}���A�n�R�V��!�>nY?�����J焸)�s��x�&��똾�n5��������E��k��7a�����'�����/�뉖�H���7y���	��ߓ�`Ԛ!�A�K ��HsE#�������d�{,+'�:x_��_kz8��e� �{-<"=	�9e+�l-s��@⮦�{������v �E�Zg�����(+)*��'�ǉ�����M�`��J��j���n@����Q{}���@.OĀ�����2Q���jE�q��;��[��'����-���H� YAA��0?��h�(�Ȣ�Q��7�j�Ş���G�(�:Q^�W�tyN��tI����\Դ�Z��0"��ZdR&��"�a��I��%�
��
�d��W���0.�2HJ�7�z̊�v�\#�/��)��T��}��	��G��9y`4�i�MPϝO;'y�=������S_��{�VFQx�)��i�0�jF߷��*�5��8��wduY&B{#���>�w�dc�B�_�2��~Q��h$4q(��iB�S�.��HD��T��č�����aXL�B����֧br�쟹R���Dp���O��q�(�Q?nrk��zO�#zd�;51�?��/9'��K !������蛠f��_goJ���o蝸i�HSJx��oX��V���BԦ���n�n��Dr\�C�U�=���3�G�z����ݮs�,��f3��V��b<0Q�` R���v� Q�*:g�����7D����&+��v9���8�B��ǲQ�����e�#���⃰���w~yc�DɝG�����I&��ԍ�37 f��P���'A��?��>Y�����l�=�0)|�X�zw����MV޹x�}s_���NP�xOAOoB��Ȟ�瀯MgF�?�J?գ4M�#��l(j��*5�9�*��uZ�R8��]��i'��B���ȌxC�I-��pAi A �}��p�^/��`y��B���T�|Y/���[hS��/��?4ެ��L�bsWQش/�1�7�_k�
�G�SE��T�m bJ@�MH�?�`�'����%E>�v܄G*W��!y�}�,��o(��J H�f��įŮ���d�Zؼ��Z� �ǎR1l'�
z0E���l�U������g9T(�w�r�^�����`C��m���O�QN5ŷC�隠�$x�ld�4ސ�@��^�C�aeqMZJ����Bed���~�\�I�Foi�S@F���t�yi���)BG�z�B��//c��6�,Ti��|�c?6�kX�Q24�f��kWIਃ�	\g�h�=�
6]3P���'._*��e�*-8U/��c :t�S����R�
WB����=ɭ/����A�i ������{��!x�C�4*1n2Jx��K�Mp�/+�u��R��%G���*٨;ٳgok�-]�=b9�#^�+Z ��G`��\P�z�Ğ�F�rvN�V�\���3[�m~�z�ʴ����A҇�R4vۘZ���X)�[�**�-�^�^]�ٺRf��z�d�B^D[2;��&�O�]C4����2��(�C������x!�ck�����[���ӧ��fӨ
@Y�C��RS�9��q�V����Ѭ��n�n&��Y[P�P�A8��y��F�) �I�ֳpȣ�䥶F�F֟��=D�8���J?��
 �{i[L#��3�r�m9gv�&RK']�☱��q�5�dۓ%l�k6j���Iޑm�p��,]�6W�Ƕ�����NJ��|��G��e��]���GO �_+�r�Nت�j/����#�f5=��o�g]|�h��6&��"��H[��Vž�k:smgdgVV����~ͼ%�ڂ+Q�g��W�#�X���� P�t��a��|��/3S=��4ڣŽnh�ʾF�~=��{ݵ�UU���F������s��x���O��K�p̅�Iࠏ�Xv�k�0i���3v�8Q�55��g:�Ha��V&^���#���={�S�G&�[J� �H�h���"bd������y����݊�.�9&�D]�R�Y�_F�=kr>T=g�|N4a:P�~Q,���sm>��0���roFMj��	�ݢY
oy��\��Jy��(���N/�aN��A��[&���N#&�lZR�r�	1���^/��O���0���_������W�v ��W� �m�G8��äBI�Fo7��B�ê.�83�	Q�
����r�h%{���=>ת1�l��a4�9̀?���P��p/,2t��i�׬�W����%�j0[�*��{3E^�������6����
�ڜ�^�cv������~�;��y?*1x��-�y*�����Gu��C���D���xw�s����.��xeO~�����e+txG�\=ڷ�ǭ�'^�E��Z���o���,��B#�>��s�hqȳB}�;���!��$�j��l�U��	���?��ln����&V����NTYa^ݜ��5��1�;�u�Q0��X[�8s��g�0�~�f�V$>D;��E�%��$�륦�4����w�����<ۢ�̈́M����K��fw�Y��Qp������#<��be����1���s�v��X�B�B>6���g{��01o ��88q�B��|��\�_Y�||fI{��.�(V�O�:x�
α;>��X,�(�-��� ��z4)��sm=J� �x3��@��`F ����J���K�I,<\Y�%뗷N ���B�d�|��
��L�,��as/��٨^���Ct��0�d05�8��ދ� �Y��Fs�Qw�Ҋ№,|�9��$-B[����;qwx��n{�Z�O����*Ú��s!��tc3���k���^����,8M�zJT|�HDĮ)������) ���VX�m����*b�1��W!<?a���.:�Ef���r�%�x�}*|��t{��4��������uh��sU�X���\���w��u��������_ $�4�\ղ�KO՗���~Lfc�փ�mggNu���y��2��C�~�:	��x��+�dΡ'gi���g���j��&#�.����]�V T��������'4�:2le�$H�u��#�e���w�&�'ĦPԑ�MT�fO3E����qY�X!�Y�DF" .6<}R�FdX^��ױ�T���+ �o���02�F�Y��0�be_u,�ˠ�ˢ_Y�[�i�0�'�+֍)@=T�]��$����Ō�t������2ް���IWhP훋2+st����#���8msy�ˇ�y,p%��� q�~+���V�J0�?��i�*�:��t�����!��Yh���Y��0�??��Ĩ�8�G�N��'L�%�X�>����]�C�
�tn�ʘZE�a	��0mѮ{nD5,Ov��΃�k�f��9��h.JY��I���.�F�����0:��U�~���Ur��cI���-3�eVQ�b��0��1y���Wf?"���K\���i�����w>5b���������zw���7�'V[��AȀ��%�GD`d�&���[!��~W�hVqc�D���*?R��*=�����}hֽ�SK!.�m��S����[�:~�]"��A���n6��z�D |uc�m���vC���;.q�0��L=	7J�"����P���QR 4��}�uݛ%��;�+����"K������f��f-�L9Z���l����bI�^d�;���w��w����;����KȾhf�4��W�%�� \�����m���y�Z����Q���>��}�i[c2EI���u:���ŝ|�𳒆�<US1�*�փ��7[�r��Yb���q�|Ш�i%|�gFԮ������}�\I�WE����H�����'�[�+��D(e�.�A�(�[��!$�fͩe#dy�w��k��`c���x+�3��:ݰ����b�*�>�`��l��1sD�����z�f���"�R+I��"��w�l�K�Dh(�#L�w|��R}n����d��_{n���X�A�	�f��?�1�(RR����]Wu?Zb�!h�7�UO�������Ec�7�y�p��>���0���k���+s���������%�όl�Lu�����!��66~�<��a�tt�ɝ��P�&�0���E ���
��n��P�h�S������V,�?���Ϡ|�V�
�?SN*�G�8ְ���L����6��bWZ5�Go��J}�3���u5l���ë�z�ym����G�M�Ov�"z�[ Kr#�qkD3:5�V/4l�H)�u�Zu�o1ղO+J)��I��刜���x�q�c�M�s��7���b�lbR�%�����yƼ�C٫vѼ'�u�O\�D*c�/4�C��%/U=Y�,���0	��}v�q�kl�	�	�`���7�'9pě��G�A�y{?ja��o���p=R��HڕG��+�oU��k�`��&ug���QZ�Z��"r�942��b╰�6��Oá8�;H$���i$n`f�U��zk͖	w�61�E=���u@]v!�(�:�ڙ9S6;�.�m��C�{�)o4�PB�E�g�:c����<��P��t��1E0�I����d#��0RRDȝ�]�����lnTgX����NԎ��ƦD�����^K��Qv�����r�Ҋڰ�@�7�W3������1�
�׳�T���,]-���nf왴�?��I�t��羫S���5�C�fI����8�ד��(�Y4�D�(
�{��z�b�e��&&�л-�pE����+h�hFU�ŉ���}[�C~�O�Ԧg� U��0-jd,
�(�R6y�t�c�`�H��˔�I�M+p ���G�M�A�Գ�W�v��e�x�Ȟ���>vwU�����[��2(�OcZD`�[�[](�1ӽ`歋���W�4�z�_�خ8����5ͲZ��k�!�M��=ጄ�,�Ah?���w����k`�@�?.��%1���P�����Q9�1?��]H�PQ���
�ۄO2�&@fn����*ؕ�Ac���u�]��0oD�{s�p���婚SqÝcK���jx/�c�Ř�2�gޤ[���ae����fhY��q���y�W��:A\*��5 �Q#L� �Bϗ����㪢�cL�P1ea$��깥0�����0�>�;�a!�;�����G�VN�T21o>�mCs��"v*��-_S��KVO���w�3���,�����"S����~�h��=+����Z��:�14"��(!�Lf�+1.l!W�w��$���W��Q����K����6�4�_�x�u�̡䁯(�[jC��G�j���%��u���9��BʝY����"y��A��zJ�_��SI�����~>7����H9��_�� �{(�������7[�MZO�r�v.���DV5se�V�<>�#�)�E����S���<�����rVR-���E�]��A��s]�ӛ��������wW��hf�;�RC����4]�(i��S�r>� UN������H�U�o�
�-�B�r� �����{7�e�TW��zR��Y#��<9k��9i �x�r���0�k�U�/�.Nd"�Y���U `x�t>@6_��D�É�l�B��IA���>����A����	��CZ�&UdҢ�C[��<�g��{3�[�9}�����[W���"Cj�����������]��φ�;�m�J$��{�F+O?�a�'�= \t���=!y�j�ۻ��? 7�L�}���K$
 ��Va��݈���`"��#��I��!+�+/ �P�\�	��غ���� t�������.$���9c�!�	��I�ᯛg~�Mg�:N��A���R`���=Gy@[KXt�1���e]���1Ȥ��ˤ��U$9t:��/�O���� ��V,��gSUo�ANd7ͭtO˚D�	�r&�o3Xr���Y/����q�}�ψ̖/�3��jB�@hI��*u����O������i�.1l"p�f���lL}��[�\�����5A/Vx���髝��f��­�x�|���l�}s3��պ�~M�m�6D�U��6�'���p���=FR{�W����q��H�����'���oK}�%鷈�&4��f*�ϖ���2���,��s��(y��ld��St�P5��#G-�ϟ$.}j\#Q���C;'��PlB�(1�0W��������j�Ei�M�������AX'�LȯC�OD�Y�C�Wcfs�r��7��^�c��1�3�R��*H����z�.�>?�,���+K���i�4���ӊx�bB*%�������vYH�g �e.a>"0�Q�V���H�L����"��JL����j`SV1�V�<%�c�B�h��_��=��� u[�-���tlcڭF��F�`J��
��eGe�(hK�0�M�T�Y�W�T�qc.�V���"�,o���B���F�[���6]	*S���-��v D�+���(�Շ��c�l�J�m�O�7���u߲��e��F��*�P����0��k�0�����=	����[W��'],QV�G��W�Q��?� T��=/{�-)�y��t�l\Z7c�Ş�c�I9�Z P;�$&�Df2�o�c�J�������ڰccn��`+�ymv� b��g���M@��{�*d-���.9G�F�P� ��~	��^�Й���y'E�S���L�n&2_�
�/����o�'��e_��(����ךm�ڄ�ei��:�ҡ�fi��ZCn@ cI�7~m:���$eӟ��x�;u����R �s 6v�>�Sӡ %��b�α;sɿH��D�^�|:3ZȺ���
� 䤭��Kh�v#�S�cСb�*�'�Z;����qq�	�'��J���\��S���+�DK�;w\sZؑ���
����HB,���g��P�=���6h�K��F��5���h%�	��Nŧ��B)� ^#,��1��,S�� ��w�,�`��E����
h9L������cB�@̆�ꈌ+d��t�k5X��8'�<���N�R������A�F����Ӻ!����5Йc9�:I����@�6�Y<�Dz��WL�{�!_Ҹ��	�}h���0nanS��%�˹�f�vb��)JE��@���óv��{���5{)z�;7�$�O%�_c/�x���\���&�0��ʃ?�ig��#<���x1D��C�s☨��
9�"���:����@0 �i(�ulJAX�cM.^�r� |�$��d�F�l�'h�����
{Cy6�1��y��n�zc>�; �N�D�e�gՕ����W�c�i���DuF\�x�80��F�:]c����L�y m���o�"�c��*�7�@��P�	� ��[f����)�}rH}��/S���vA��X�q��5������F�eƑӎN(N�lS�<ɾu�7ѿޟ:��9F��&îս�.Rt��3�Z��ڥ�m�### GWR5�6%u*-D`�����e��~��Ff�i8�ow�s�6���8*�Ri�4<'i�����L�gpc��{�J��	��G+][p��D!�C���~��K���4e���y���az�׫���3��v���3v=4�7kzv]8َl��(O��Ib>���R��E����-T�>���3o��d��pI�+�Z)q�"���@�U�t�;T�w�t�ƹ��"QO�
����)�X+Q�u��.u�Iu��׃��U�<yY�>�s�!����w�t��l;4Eܼ�փ9�|���4�{s	��AJq�(�%UOp��R�HCl�e��`��zA���=(�x��l7Q�93��ʢ f�erc��y��&ƾ��%b��E>� PjJ����v�����|�	���[Ӊ��%.v��1����[�+߼[�e���"-0��O��Q_|�Kp	<�g�)��y��x��Z5��������7�Z���hi�!�
��縆�`�
�Z�]m�}~�fK�a�7��$3���%D����B3!�� ��W�	n�,���P9�*��#谠��`Z9�fE�t�k�H���0�Z߿��*!��q�=����y�Xeb�HI;��,kWÙ��G��a't@!��B�V�i#�׉+��m�L�p�!��E��z+�����&f��l0���b+}��j�~�}<^�ZX������2!�,���D�4�r@eB�L)�Z}��&����z���1V��5_6Sc6�#H����8�$���̚�$�k��͋7�m��˒�\Y-�-o/{o�y4��
�t�д@��I
�\3�`�(�����ۈ�%A)̸����>{�n\lN�� ���+6����e��*��-,����i�0���ke�^,���んѲ��-&sEon[�>���g�X��D�\b/�
��p�� �f+���d����9O�4�/j��B�/dT�=����$w�
�Δ)�
��g��I�,;�P�Ǣ<��
�ڷv��9�^��҈�51r@�����ʲ8�$�X�J�LND�#���\��+�5��hj�m��	�yy�4]qג������r:����.�h����N�K���%�rUV�Q��|*ML֑�$}N��=+}��cP� ��5�4�0�5����9,�
gZQ�&Q��?�J��F�����.�Gu-u�P'�;��S�l����>r��8���7�;�(!��,��t�1-&���h,F�6<+z��ʽ�#c�E�5�[v�܂����r*H/Aw%u�tM�q~`~����
��6-6)=�o۟���{�[����]�z�����@aw��-���v���aW�-�c9�q�
����?w����j�r��eIsӾ�"��0}�V���Hs���)��d#߻O��a�P�C+�"�o�Q #F �M�7�JI�	�-��B���eI�9�c�e����	�!�X:����o3�Ac$k1���H�B�A��2F75�Ύ{��:�B���&�$K��b�E���jˌ!�Zޱ˝��Z��[EVU��")n��FeO,X��$O��9����]�{���X᳊��<���z�I��X��Hր��.Q	7�'�ǈ��6(�@ck��K�����K�O̩�O��QO.���O#���gӈ$}cuP��&:o��4�W��9Fk����a���f�)��d,LF~x�L����8�t�K��6W�P(��6R�1$e'�����G��|@f�a��|U����K���S�lL��>|��ݘ~��� ���}��{�y�H$�.�̗Ury��� �в6uћ]ָN����_��(�g0?�;�佽�d$� ��p��:F���\�#�r���jW�̟�3�a|���+/p�\����#�J"�DU��x6����$��>uO���lӽmS���#)���uƳ-��������>�G�� :z���w39�,���a��0� ��%ӓ.�'�J(���F�9��}F����BX�kG����C�şh�o�����7�2�e^��';ׅ�7!��tm�����F�ބJ%���*���Nؖ$�v7pzt?y"}�1��X5�v�Q�yL]��
�4�!�Pd�Bz�����X�&"ћ\�mZ�;n4�BO�?) ��~���c� "!*����� ����̪��*���gfE����8�\�H�������SM
������W�w�cе�_��F���)�`Ͽ8���;E1Z_e8W�*%����"�8=I�,"q-�H�1��,�h�_;A'��`��7kc��P�]����<�i:��E$@���� ��]F2����s��%�O�u�5w�!�Zr���)}ݐ|e7�&����o��!ڣs�r��t@N��$a���n�^�wc 6
s���̓�O��@�:p��@�?r��$�}����[�#oP��۫/��G�����ᙿ5�ĉ��<a��+tq��y6P�y��C�ܻ�s��f¾�u2��"�FX�{���ǝ�t��&*#Rȅ��&�f��b>���x�|z�7"٧���n|�����wz�Y��<�Q[h	\��發���L�|�� �(H�o�k�cp��/�i��J���bV���z�PK28����&юE��OkV��A�mE����Gj]��sw�dK��_\�f��\�E�h�nC
͆ԍ�E�>VA� o$|���(^D�Q=��rfWf��=������i��rhے�.�	�����b�)Q����)60$A���h-Kj>�{J(`P�gg�۳�]|����4J��v{�0_(���Ҷ���2a	�$� ��Q��У��"Y�j�*;�0p,j����p�
-H���iX�����#��XE�Ļ�[��O��zњ_�P�=V��_y)Z��1DL�B��®�[���d�q�sj��-�io�\nn�,��\�o�m�w'`�IJ�p9-,�4 ���G�l��ǯ��+2e+`�e�{q��@S�vS�tɰ�IR��:��˴%b:�u%>�g$��[���D�y9 ����?�fBV���n2�>*�4Rc��Z/(��V���s�N_�c��Z����dB*I�$ ]ZkE��]��@keB>H^j8+�4�N�ϒ�������&��*<k��
Bt�KЫ��(����R>�;	�u�}wǗE��$Ln�VN5��ED�Y���!#"Ujw�m��c��� ��M�����ke�#��b����9�;��MY�;��(.^L}�<�� K�n�|>�h��UEfD��>��Pߕ�Z�щ�4���"��� 8my�_�o��
w��щPJ���]OE��������i��хm�K�}��+�������/�=�g�좕�lvԿ@�K�I��O���;�qy��h�uW��Y��z��صMc��E��5���#��3�ؓ���s��=-t�X�#��T��=�N	O.�C}�K������蚏�qc�\��]� a!�qً��Y9t{���'�h��������ю�w�4����7_VapPJ�O�^�HEc�9�R����WB8H�B͸�Ag�a��]d膲���2��({~�e��H��PU�]*�\�g���y[Ӧ��!�#&��.�D��f�7*��%�R��s�(G�'�f��Ѹ?E��~�����Fu���ܖ��
���!�=�W-7��Ϊ��E�4�R�]f*!�!���q�l�ilr
,�C�1�8�C[O����M�Νj�ل�љUr�nk{��Vy���D:��U:�z�}�{$o��'���P��x+���sn��b���b�M#4 ��Z�c�)����]4l[-4��s�p�PI����J�lRhD*�Ɉ�f@�[V)xRK��جs'��,:.,mҢ6�C��s�_��u�d'M�՜J1j��g�ZAd��q#����{i�~�����rÖ�| �!d! K�A��?��/3x���K�7�Y�����n��OKy#��� +�k���P!��Q)]D.��3e8�r8����5%4���I���vl ��+�vϹ���K��۵w6	]�x����h%b{�m>��M�oi��;�5\�U��q��ϙ�Wt�.�6��/M��n��O����?L�m�TbN�{�:7Åv���������7c�ׯ��l/F���ы��O���V�ګ(��G�)�~`��\X��H��#qoSn ���Dug|�(�:u�`#����,u��sV�L9Ep6ؕ�ّ8,U� �B0� I�ރnAk��[b��N=%a6�߼0F|7� �&7�
�ݦ`�v��?������w3��2��[��	C�C9��� ܮED�w�P�l���7;� �n�'g�';���9�)��� E�N/d��|˂!'�1����;�n7��D�r�M�g�p�>���a���L�K"��F�푾�U�T�v{�=�4���}�7��s/�?��;�;��4�%���'X?���/�9a*���� 4��8@�]:#���
9���n�LS��PQ�i����c��d:וF�HGm�@�&��!�V�T�m��`�`�j3(8�$�d)Us�6����=�n��0��ތ,
�b=L������i\7�?�@9����&`�^�E/�dG�fw���������x:Y��z:Ŀ���^���D#��	��w�kR���G(���kmf�t�3@�q�R�R�.��&0'mq�t�=j����~U���8)�R�o[gP=���Nk����2Q�£���4C
ܶ�ӡ$m�\��m�!|Mx�iNV�i�cGZ��;��	��f�.V�d� n���!p/2���T��X��I�M֠�+��$g�PTUn��M��-bG�R¾f��o;y���94i:��n�?c�}l����C����b��\%�cU8pP�[�Ҁi A��ԃ���Uw�>���l���c����G�h:$�����Ϙ0��ЃRI)�U����O��Vܖq�Ю'AD�{��#���ymv�	K:�ū4.���	�S��hé�E켎���a�B�gi�������x�dIސ������R�T���H'٩�U��y,��vC�-AH��`����d�2;O5�2��]gw�Z1�&?Np��Z��G��	
�������x﹠}
j0Cځ�PI��7��*�G�;�{l�4��+�r<�=�p��oI��l균֮Fܜ�1[#��F%)�%�����=nA���#;�Ȋ����>�l���s;,�4�~��tS�t��a�Ϡ@�>m��.4�Cn�
��Yvx�c����6��/�x	�WX	'�@f�`p@�2:4n�AP1-�O�}�:��P���U�#J�G���E:�,�Z�S�'�.�a�XU�dW�y�h\Eq�i'/���[G���m�������+���m�~�YI^���Ŷ��l��ץ���$u���=����㫕��nd�Î�Ó��n3������0�1Y��)쥍���s�ڽ�����ʱ
L���N*��G���'|��f_S�c}@ŏ�Cb���l\�?W�Υ��e0g3w��� ��=#D�!I'��6�_�u#���GZ�Éj��x眞�e���� Z�i���̯����87�.�ZGvvlh2'�Ξl�O`�O�����͈���n@x�s�+"������F�==�޽��%�Y\��WQ�nP��n�22�&�� ;��/ܔE�P�LZ�Wa�T���S�F�s2����Eֵw��ï :��y�G�%�`y�N5��fe !6�g��Pp��qb���Ck���ST`�� 	@'�O*��-�-5�{��	Ƀ�۔�gd�j����1��"�J~�Пdz���=��o[�E�2�C~m��N&*վ�lż��{6v�~�^��1gI�Ŵ���F#����&��hmy�xL)&���҆��V�\f%d��G����*���9{�ǹ�?�{�L\�?�� �LG�|CO&�t�(�1?�2��C�2���c�E��G,_��x��1�`U~����S����<���$��z���H��r��j�����3�VnrZ�$-z�3ߌ�;o���o�UDCs���zc��B��1�}�lZrŌ���ؿ�2��#��cj��1�-̥z�
:���c�N���aI�Ag4N����������s����뺴d��� �m�y����U0�����K	��m��C[��6� Fj�����^����wo��ꓐ���57:�ZJ�qe漼J��ή���M��a�ܠ�/Kn"D�<z�/�}wk���ru�!SFy8Jr]��F)���E����N��]���9���P��)�ˈY`��{=����Y�DG�`}&��0Д�ט�w��i�~�{f�j���7��iJN)b�S��H�������ݸGB��DH�Ei�mv ����@��3�U
n�%]�J��U�b�o��b��HT��Z�nYНJ��s��|�.�h��&d�.K���x������3��$�'�Q��}%��#-7l���Y�o~�i��a�[���S�q����2��l}��(�k|ڟB��D-����7���'D0	wx76�⸉��O7L�b�׳uъ�OtMimNV��-:��-E��N=�LU�n8�׻�y҃�kp�s��|M���MJ=WO,���:��՘�Xr�|�O�Q�75�Lz�����_')@���6����O�OIF�"�/�$��iǖ�.�l}�@F�����J�T�}�)H�S��ˉ"�B-(cW���<ɫ�Qw2�kڂ=.�B���.�^�w�D����80ih�)�	J�z�A�/Yz�yiOctd)sx�d�hL�[����EptĪ����K��?�iuUD,�h�@���N3y� a 9�W���%X�P���H%O��>"�i$=���b�c�u����]��;U0�c�{����T��;�y��V�'D����ˢ���a-�����ݖ�a~&�z��h�-�~��2 �tx^�Z�w��<�u����y: �|��"����
�>$�T��$����d~��tz��dK2�x����А���G��a�,����Qpp��h:~�%[����	�Iڔ��ӈB7n��>�m���v�����H��o(rb<�?C�|��K�#�U,�Ɵ#�#�Π�nt3v��?)O�nWO�������yn����m-	+::9¹x�^�����..	2�ܙ�gA�z;����+���Kb��}hm�K��p�/�X�ĚCR��a0@��������x�I��&��Њ�@4R��gQ�S1 ����4#�G6e��p�c1��_E��6�9�=0��l��2��su��L;G�Db,_F�d��?&K R��I�V�K�Aө�U�2󯦻@��d�����]���� 
aT/��@"�tAb��R	Dp��0��bLA���fB��b]K��߯CHH[S!��I����5��!8�K��u�, �d�{�<�[G�-��u�7�k����	��Gw� 9�e1��m�i��������6�F�3�s�yzą�a(fȋ]��GB���X�I�1=��٠�q�U�# >�P��;�����ݍz�#j���Hɿ��Ov��Е�yw!w%�c�A�����Y0���E��6���#]ko=�%��TQ,m9r�r͙�d���JN<)"����'f���B"Χ�{d���7�qa������4/lL���)�i�LֿE�L��(����>���g���|-aǦq����h�$*\i���|Y�%Zu���B�V�8tg,��:����.;$���!z���nƍ%���A!�Tnp�)dק��2��:\��a���`�Q���=���SE���
/�ʤ/U.}����Bof�_@�vO1 *2K@�42���Ŧ!岉@d�C�I���ݢ�|~ͷՒŰ=0�KM��� <%�W�U�Ni�ʕ	R�Yb�z7���ˢ��c�)"+�Z�(�B�Q�����\x�*U��d���N\+�X�·nt�]Y�kFʮNa�����o���Q�x�$A缽����� ~;�x�<�gC<*/xA��6N
}H��>b����x����U�町�Yy�1��X��Q}<�b��LPe�- �ȏ�[����Љ;�G^�����<399����xFL���. z����H*		ׂ���(��u\B\:�
y�&��hZ���Ch�h�|c��XDW�F뵿������5cWV�L�vҲSf��J��+߂��K��z�[�� �U��n���sd'�yjYU��oN���Fm`db�$$�4�+n��Z����0�ل�FJu���8���&�-w4���+�y�ǔ?�8x+YKD7�=��ch��]�Eow:�U�<GC�7��O^U]g�^�I�gй�Ӽ�ŉ�i�,���0{s��5�|��|ܡ��΍-]"{�S:aO<<�=�8��@�%T�M��Q�1Mp �U)��҈�N�ɘ`����O^� Xq�9,��p��$j�p�Ll��]}�;�߸>��s��$\�Un��z94�h~���\4���BACZghC�<�\r?.4���tGL��	!<�0�w�B��F|&�U)��<�����9a�F��XpB�tf��U�3{�A�C�\R���kS�$�N��b�\V�o�Rt@��oL��I�,���e�|�9DZ���,�pb5�RX� �����Ju�~VvH�!�X�R��1D�t)��+�*~�z���1�����W�O��� �p5�_#L���m��w?�y��$`ZkB��^�)��d���,�/��e���).�K�f�ܕl�x��쟘 MK3��k)��n�5�l`��+3{�A�Ǌ���᭬�]y�{�V�c�#zڳ�V� ΗhJM'�	?q��=*�%v�?��>�Ѽ}���cR�pިϤʒ�J�729�b��d�ڨ Zو���ψxʱf'��<PQ �5�~;����R��ȱ�I6�z�����ڽ�!��SO��e6�$6)�F+�@aN�3^�ea���I5�E�h�i��g�X�/�qp�P��<�P{�1�q��Q5�װz&�	���+�bX}�W��۾�ּ̹�������$(�%i��.(��a*�l��0y���ݜY��Y �V-�(����g�k)��o���}n���%#},�D�.��C��I4)�,���� ^F�_H2��pS���1!�����n}��cW�j��h/v}�5��<��j(��'���$4��m�VG�\ѭO�_K�SĲ� �f"ȗ�򣎮Ն���`���D���W�9eN�Y���5k2�:��߳��r�u��jW�0�~�q���A\�4���1H����%+B	�8"hUR쩱�L�%���1��g���?��
��x�/Z��R-����!}|�bo���7N��5�$h	�M�<t���x�:�a�ƒ�HZ���}q�y���ut��"����k ���b9w�'C�����w��7����JZ�R�����D�dP�I
C�H�a L��4a���5��PƉ̈��_N�)���U��PB[C�b��$OV1u�<� W}���(L�B��b_����YJjr�*�[-���v�	9��jG�q{J��t�<�.8��<��$��ft>�3����y>�p'��r�<����jaE�{��H��t��|����M3F��us�x�L몐a}~��ט6�jCct )orE����_I"��a��R�v�Ih1�RjW>��]����"<B��I�(mxx�_#{�|��5q�;�"�+<�M�ZΟ�q�KH=4J�V�����a1p��c�Q��<��H��9�=7 ��Nr���W��x�{�-��ƄNZ,JS�̮��BT���Y0UΓ�ҍODڋ�M�}��g��Ɍ�İV��j����P�Q̆�#!"g휰��߅�	Ո�d��5��ک������.�IQ��'0˅
i�)���S�\G��x�?��W�P�F0
{�\�ž=�j�C	\�~��յ=+��j�V��������  �������d�#	��=}?ڰ�#0{���)C��Ʈ.?�%���^��֋� �q� \q2Օ`��Da��e�'m6�Y>$u����G��*&!UP K�D�
v�>�ۢ� �I��B�׉,��J��pZ<�Z�|�0[�O�����5�{����n'4�g=6�ՑF�Az��W]���'~rf!`!v�{�S�\��ݿK@�o.OK>}3a��>�s���^s���.�`^!�m��9x(UӺ�!���P�\8�������'w��I���Qu~�:M�h�6Z������˰���n`�5C�m�~��-^�#D���9�N`b���>V�=І������5��Θ�&0CF}ه�v�'�.Ru$�$]�㛯�9ò:��Y�Ao����A"Hm4���Z|+�F���j�7���;����b���\+��+`SgR5C�ib��%CMTW��GTp�5��2j��%�6����:-�d�2i�'���c�<��&��n9i�H���R���!6�!�"�Q� {	�GO��(�����x�[�Q����[�<�"<x]������X:�h�<��UN���,�LO���#}�n�����D��g���� ]zZ�N��E�j�0ފ�l���B���r�L�ݷ~�o�9�F�f8����:�/�?�I��!���sh����@:��}ߧ2�`O�_!�m��]7�[aP�0b�R��������i
SM�S(�iX��.0�Qs	�l�Z웮���ș���5I��]ߘIlIbUb��6[Y&�̈�>
�H1J<�n��E���Twwp�> ���?	tJ�	�$! 	ֺ��c` V��z\��6����G2�)�k}X�:gW>1�P�7�h�>yD�]���5[[��Fsc��բ��;�sOړ��F ȏ�;����N��Au�����Cj��v'>7�ԝXĤ��'P'��;\:CI7��1˩ui�1:}����]����5�l�e���Ehs/@^&��+��0�CUșA�yt&m��uǘd��P���:�ߙ�=�v}�Y��`�/�� /u�`C�?�7K·>��4�������e}��n�M���3}��NK�I��5�I��uXɪ
�G$����9�F���do-z&���UV����@��{�g1�R�x�Լl����Ok�Q�6wV<c�!.)6����>��u�;���æ4	�����!�n�4ba1���&����ٍ:_���s��M{O*9��D�&z��nL<7�j(�	�kP�
�d�8S�h�.T�_n�I��#���HW_�'J8�O�J���3wN�>,D���m����XtI��9���.UU��.\���VD_���[
���`Bvm��t��R�	=��.��Mb��n�P�_lo%�>Q�_uA��j[A�_%[}��Y��ۃ�L@����Kk�;t+��������GM�q�_oy1?�*������P�!�wl������_גƼ���̭g\�T�`��	Q��=V��Hw���[^�g��L���5ڑ���"6�V�Si�_8X����B��Q�T�ɴa� �je�j�t���t�~kk~5Mw����,�E"�(��HQ�Ԭ����V�}x�!��˽;��8��&Q�rO-A[u�q9���=@��P�'��F��5����E��u$ kcs�h��@�C�<���dB
�0&������8�9�~tl���lE�,�����>�>� J�t��DO�	��ʩ�}j�~�4#�/��
�yp�Mm�MI.�ǥ �cUL����n%e*�1I�6(5�y%l�ԣ��.�d�R�O��O;i�������������4��z�F��C�^�S�H}<�,0����C�~[o�<�13r�������r��@��H��G�ZN8��j�.4�Ց��%ǒ��#���,G�fvy_�|*�,��Pp�8aA���6Av �T�TZ��\e�9T����k^r0彀�Zx�hX�.)+�)�
��<FiW�"�<�
�9�$N~�����@�<G�иڏ��`�����ۧ��#Hh�Ֆ46�@Q����m�E,��CMOl�G���j�'�0OϿq.�eK��{�bW�E�+,I�3s�0�S��0I�˼8��f*�G=+F{:˵; 2����1'�j	4Y�첰�-��
���8� �	R�x�VX�Z?���a��q �$���P�;ea�}G%�b�l"t���z{�i�p�ځSB1Ddʧ��iF�}�>M�uu��lTc�Ũ��MS�O&�����ڀ�n�ir(!���%�4l��t�~�B�(Mi���<��Dz�*f5ƚ!IQ�u��L��HE+�(���F��P8�e�&�D�t��"�1`��
gJ"u�§c���>��ǒf.��\�6�"T�f�H��܆�$#���J7O�>���.S����C�n�n�r:�J�Mɓ.%nH����4%(�W������J/�U �,8��bt+ab�M ���9|F;	޻�߽��%w�>h6�SC��
�i�2[�[�E���y�O��<��M�@<T�{���P�0y��������=�Y��vN|���	-
����!�4#�c��=�k.�4le�D�:��A�H�1��yY4�4�u��M'A�����&j��P�j�z������48�-���^iA�{Gҁ�з��w�/-J��\�_H�Z9�&��Uą��