��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su˸Y��'��d�Ay~�`�i���o3 1&����1\T�����	��!mF��
��\�ݘ�#X4|'�~a	N�1�""rϗ��?���ݝ��^��lt����d�k>O@�0�#/�����"WYj����i� �N�7A!�@<e�]ң�;��5D�監p�.� ^+��Rk0;Õ\z�7PF���p�e��	��j�kdD/���1M���(���T�e+qr)zD���FWkV��������\���mk�*
`�R���	j�' �� m�cD���9:�DhT]�����۶�����i����ޙ%��d7ܷ��	�:���U��(�����#���wv�pFc�o�m?���<�δ�7P����( ��(�����1���o.O����BE�l�pSX�m����
'j�ߑ?�a\����3!����� �@��+�9��d�RXG�w���=�"�c�Q��j���)��v|t8��lB�Rv�g���3���hkU��q+��KC��L�-:��|eiֈnö�ut�c��OX��M��M[�lc�z�	Cp c��~]��T���H����1cPa%��<�Vη��p]|���Do0бb,�cy���;��U��|�I��F�x.�ߒf�z��%>aP�g��3T���cU�=��}��J�/s�Ȱm48�3>Z������~�Jѓq��X1#��ty��n"��9rxu��(�4&m�V:�V�$ym"�<`�-	%�Y�`g���	���s�2��{w��ѓG�q����Ă��?�bQ��'쫖���}�k��T��{f�e���	\�c!�("�:7�"�;�
/6�冠��)"!o�g�˥�C�7&w/��،���z
c8��U��y��T��}`�_mdq�ۆs�J|��=�Vъs_qa5Wu�2v�>B��#k���[��o=�X�u� ��RT��̙̱����rH�o�+5E�j)d�Q�Ī�lGa����>w�P��mnm���o8e� ���N����z�7�sci6;�9�Θ�Q�c %��c�C<��H���&FQ����uY�Wx�R"�5�M_MW�uI/&�a���U�0��\�1��ʻ���c�0�cP�����?ld��-�3��9�Ʋ`��;.��'!�'ڥb.�`�of{4����On�����ޔ���#������ј^:>)>)ٿ38/_'-�����{��1����V��پ&���D�^P�zd�Z��\U>�N�{j!�O��ld���Ӷ�(]��۳��m�S\P�ȶǸ�^�/K}M�󠝡�!��Ȼ%�Vua���9���+AuN&#��Z����T1X./�������ĸ8�b�E���W6?N�X��lnc&7!g��m�F��B�~��E����@�[���ɜL��ꂆ�;z�׵h�ٌ¡"���Yh�$o��`�j�8����)P�;�Mh*ͣ�6���	)��D1��n#�!�T��7�|���X����P�� ���� ��, $�� �:��f�| �\���y��6X�Kw�&���b��^�;�=���������k�1�"]>>BxRI{�A�mC��cm�e���Ѷ������BP���@tg�`���Hw���,�xU�D��>97'Mo\}�~Z�[���?����ϋv��$�^D���5��T瓦��C�Ŀ�N�*��:���b%��}��h3ڡgI�*��<o�u�~��sd��?69�e.E� ������4�E썶��Kc<묎q,.�̕�A�?�fg�'T�2�F[������	���]ؤ��>�_Y4$��?3�|Gr�M����m0����d�L��x������u��=]��`ȣaL�Ɠe��5s�q�0G{^��Ea��K櫹df��$h³e���Dށ�, "��H3h͝��s���}��� ���T����b9�mQ �2�9�@��V�ɶ/c#����k����u�ε��<ߝ{b��ǎ�ۤ����g���1�݁�uo������T�6�X�5"�Vtt�+�k���ut�_����Y��!k������Y��N�6 ����d�G�UPPe�WG����
�����<B@�e�j-ɓF�m�զc�r���;^�)��ߪ���,�H�x���P�,��� �Un���s��<���-:��G*�
� ^��.C�]q�����y���59S�܁	�m�=;٧|��P�j�1b�Z��<ߔ���H��]�pP��8:���(Q�lb(��Z^�!��]����w��$�?O,�yS�?j#�5'9m�ݲw�B�>����b�޵�,�z�����Md��B�j,�cV�Jz�4�囿O4A4<(QR|yu*�@���E���Ip5�q~J��Q�'4+|�\���<HV��< R�4�ꀔ�\Y����\�LՁ)I�2�;i��<��Uh�.Q�Q���1z�%�������^_:B��p����4�2t�c(��9��FLX� ����*��J �搅��|!lg��ߣS��|:��P�J��hj�ʍp����%"�ϣ�:ƃi��/�x~�hf���|3L�̛�$Q�&!�?�JB�%���i�%����p���|l*9g� �V�<���
h��n�L�_>5(ƣ���a0f��� 3c�/�<��-��v���W ,�1���X������,%(�}��H$G&��h�֏}�9�;�q�ߐ��&�{��hLy�#�ؗE(�'��Ĺ�}DԲ���R�ri�MP��l\�	�Jr�N�kT�^f7���oL��)*;������H ��Tl���H#r�Y�$S���Z�[~���N��S��"���19��Mb�o�D�L�aE�n�b��%d�?��mk��O���o�C�,��3b�]JX�{�=m���[,��\::��;�"I{9���l����"H�1�"|,G*�Q>�(��`ص%�OX��.�������L��f���4�A�s�Ƒ
�6����~�Ռ��!��eD���PuW�n6��4�Ob!U�|�m߼(/[�yZf��M@24H��/3� �A�l��
�j^���+u�xI���?��)j���G�щ��hY�@#�Q �w�!���GU���F�C���x!��ȉ����{@�͑�<���za�S��j�5&=�at��V��dܭ
� :Q���>I&�6bn�y��#Y���^U�!�Tv��y����[������JϽ���v�����vS5Z=���7[iCt��҇�����
P�SB�^B �Sdok��YC�� �A�-P��l��\p������5G
������+qC��k���'ʓ�ί�����i,9���u0vd7�)�QIŻ���E|�W
��a��s��	�O5�CzN����6�ԗ�TK�;��j�?�`a�l�!]S�ǀ=���JEׯa��F�8�
�uJ��� �w��*%k�
��U;��L�����#��ٲ���(O>ષ����������䐒���Y�#�l�rvN :��n�P��%�?�t1�G�Q��S����^It8-#a�H>��7�o��4��9��&'
n]6�`6fs^;/J�٤㣢�# ��<J�#����Z^t��܈J��/����51��y>�}+�	�p�䋍ɢ��
9��=21��=ϔ?�&��̲2�E���9㼶���͆�!��v��Cr_�b����V���-.� 񏸍_�u3���v�.OTM�Fh�[�)�}��\+�-EyY�J�v���co�m�x.�bʗ��J	�4z�Qx���/U��[>
r��x4��Y�ˁ
�$j�|}У�Lɩ�$lL� 1p���:gFK�W�3�{P"��q%\c��ub�xD``*�v�Ӹ
9K�^5��R��bw������r����"�}6CU�,Q+�Z��R��\	�_Lˌ� ���0M�����������AU#+!���E�m�\�A������O�H���A�X�T�og�!�A�?L���a<쾒b�Ѭw#)�5��)1�G%$�6��Rq�����|
Мd������g�䶲����a����|n���V�9�VKBJ�4�F���6���wk���71\o�3SD;
��vu2e"��yK�C�w��,�!H�.�.]5�h�.%&,1��Y��c���Ne��ɪJ��`��@�R+i�Dͫ�0�����s�P8#6�&ݺ�d<6W�&��Ӛ��bC���N�Gb,�;B�r��ʒ�"�O��2��Bl�;��,d=��A���4A^"�s��S̉(����+�Չ���I�0I�g����q�OZ;=��(O1P��x&ԩM�l�6�.���@�l�W���􏰐L� ���W�K-u�(I����lCTE��Cq�)1� f�%k�eTs���K�KZ�)oU9�� ox�8��t�&�;=�7�� �O�ɩNY�#��b��ݐ�န&k��)�U���36o�S�1��{_	a�pr�V7*��֖�>B|�kuh�����m��փ�Z�*��Jvנ�G������GP��f01G�?���o}!`�4]�vj#�>4���D9+=dH����Ȕĉ�8�˸(��"��9,���)�!@X�Z�;�7����*������SN��;���V4��K��/{��j��)�1��Ƴ�7�\b�UǓ �mv�Љ�4c ��0/���.��>���(��_���c2��A�*��y�ݎ4q�a�䢩����h���I��jv-~�$�ؖVB�㛍�}x����z������l�	�]?vN��s7��n��7G	svDX=:�S���/���Ã�4.�sgTe�y�/,0�"�Z����V�*\1�ڧ.Z���T}yN�.��b)��Ra��� ��$�zfea^NJ����r�3ܹ�#��$�u�c<W���ڔ$��ڱj8�����9��	�|�#���F��a���B�T!77�����@�ww9��/fP�3����TI�L�~C�%�$	�Q��>H̝��W?US���,���J��R��)=Լu"��SE �����Į#we�J�#';�Ox���%���v~0��r)�:ͩ��ѱ~��\KH+�?��D3%[g���ҍߧNr���]�]�q�L����m��-������a�aG_*��N_Ekc2B�Mb� ��J/.*Ia��5�^�=��f��N*��Q�ɭu��H&S����!IYq�[Ծ�>��4��P��Cn�ܐV{3)��Qtx ��s.%�����@z=���p
��0VH~#z+Xv���U�<۔�\��=��r��ع�:�����r+hW<c)\����W�~��G1I�Y0k�uM�`�>�㬷�~n�)��6p�M'���R�I�>B�ц�J6����,��Fr��U��i�'iYR�駂�Ȳ�|�̈�O�g�a1�^�p����<�[8��.�*�
�Î)of����K|VzF��s4�8)6��JK��U�d��B����/��e�H�K��V �q"�B���� w�u�"�R��<��^pe>��eݎ�C-vZl�bB�\A����{����,�F��u���v%��T���;�Rh~dsB�U-����3���s�I��a���p�&.�3O1 b�>�|�G�<�^VG ��$Qf��$-`��>A��1�@��T�Hl鰾����(10���ו��Bi���L�,�X��lI��pz.q�b��'��3>�e[7��,�玚�Ť3{�He�K��	V?XW@��p��.1�yB#�se�8�?�aTB��Р�a:�o϶�r�`nȌŮ��M��-�Rp���9!eA��o��w3D��sbJ��C�#���P<Cᬛm��å绦�3�T����+�@z&�GMD� ���!����x��417Ce*N�)�2t����h����$A�`���'�^+�]�����(\Zx��Ȣ����#@���7�y��7#���a��fqD��j��?���h#�N�9�sO|+<(����3��l���B�/�a�<��5�Ӳ�T7�����]��sD�0#�w�t�����<�����=^�e��}��u�|��{�WK�7����%]�Nu �}���P�������/Ⱥ>Nh8z�����������s!�>�j��a�%)o��D�ěH��^4���}WNx(6./�n�f~��w���U^{���im���*�O�%��f*��"�az/���� rf�����q��c*�D]l>�������@t�M]��!RK$�)�<PSi��E�Dh�@}�ܕI����s�$�
[$���!�����D�]�!�Ζ�t�?�����q���N�G	�+��È<���R7I�u�<�]�$PUj��,��:M;�7B��3&/~�,� ����<�0�F��_�ȹ�[�S:�H��� �j;���=��?�H���G�4kH�I�����G^��~�p�5St�(��&��:�21lojC���6�i�˗m]��%��>U��j�|+-��&O�
�3I4+F���d&:��!Q}�)hov�x�$�u,F�G촛�*�+C��n�X��S����^$M��BB!�u���{	����{Y%x�
堊� 
�x�X�����6:���Uv�rQS��(Ӈ8B8�^A�B/�Pg���{$A��q8� �u��������=n��rL�X�wj��9�3������6���>��<����縚H��"���π��6|���k���^�9vb��3ԋ�hu�S�_[9卻iUw�u�8��Y��d}wp)����q�s��-^T��^�t�ݤZ��D���Պ�@�Ċm;$���4��
1r�f&�ac��B����z*=�e�؆��� *���b�ߚ��̚>u�����W_{�^-����F�rw�p�a�W�{��f��MS����:8AG;[e����,HO�ze�m^% DTn�=Դ�����T��C��Z�em�dN��VB�
98kP'������ք�����4'��/y���p��Jኺ�lS��(lp}��i1~ؖb��-�dR|�@����y������[i�O��d�S����o���,�૑��bI���0��*�;vW(���O���h%�@�R�5^���R�I$���^ނ{	��{��BȌ�#����"˧Y+=�2|i�����y��G�N]�u�~�eU���*�D�c*�Ld�U�u?c��ע[
�%e�����ւj�:[F4N6�#�#���Cq���m:��0;�4NP�F�PM#�^<�B�6���O(�ŀL���.��l~��Q\D�F��N�]p+���9�<���e�R�RU*i[�O�w\Pz��J�yZ �!��&~���=��3{�g�~�р�o�≞�ϗ�ע��}|�g�ZD�!5�j���=���10��O_GN��S[��!(VλOh�\Ý��<MSĞl���L#�Y��~���U�Ƨ�9���JQ��b����y�6)ϸ��y���m�x�K戮E�7�'��U�,:qT����+���b�pd�_a���{�5��L neI�3
�bHy3
7�����N�v=xX�YVv}8��Y��;���Y�u��/7)��!2�wE�==�!���v��|���p�R�3�rYzu�ϙ�~�-�6Y�$
�qUxnb~/R畚M����i��/pJ�g�T�ަt�����D��V�ar�<ͥT=�Oa�U���� �}�5����sڑ=(���`�ר�B2w�uU��U4��0B*Wg%��'j?��B��c�sg|���a�m�2 �����4
)_(�>��z�pu��)R�~��l��8�M'�Rf���R�ۼ���u�7�m�G��p�o`�̸�K:R�Id��aSō׎Y���M�Ⱥ3�7e�w�Ѽ�'��Oau���,�):���
��a��t� '�5�e�( FM{q����c��,~���[���c���Ӣ��Y{�����t��lq�DG�i�G/G�F��	�Y*2�7�a읉X@sO�f�C��s��N��uW�[3[�{�c��Q)�����L.�Q���ⵇnT/��@���@�
�g�h�Qpb�E�#�	;�&m��e��SӃ�����1F"�Rޛ+{��Fܷ�h������|��@O�T���X��gӗ� <o=��Jx1)��л��~c���Wu�E��4N�+/]�=/�$��*��/���V�;�<�f����C���#Ԯ���*iƠ̈�,F,gIw�.�Ԋ�������0ȈX��̋�,òE��^�V��)���	s$�/������Bf#M�'��]_h�䏲w���oקQ��[�
j~�_0�#��Z�B��ʊ;fW�����ڬ�s��Ȗ#l���O��޾4��:�V�񺄴7����Oh���9w�:�4(O�Ed�ؔ�P��לY;�ƬO��)Ը�nS}N0�6�����~6'��Í%� �f�2C�� ;[�r�7�j�j��3Y������� �F�q��ۋQcP��vC3,O~��?�K�b��"��C��`A^n����
�:M�dJ&�w��r&6Abs��Vu9����sX�ۉ���JÞ
���eL7����R�tjݔuL?�xx|8���5�}fd ��B��*�Q���1H΁DP�/������ 	9����4X�z�=!�����>�=�<@�ZX��P�Z�z�7�q�颋$��������pk�QV��$~��UTv��Di�z����1�P��VI��^�G/�����5N:���� bI��O�7����V.3BL��#L�Ft�O�W�
�웢������IE��^=�*NQRz�/m���=La�M���y���y:�Rj� �̈7��%N�P����LB�<�3�LLv���a��D��'vUzԬW�켪i�9�T���Wj63�.6q�l��m5ڡ���ǰ<�E���Ue2�O�^>']��,F���ڝRcۋ��,�y�,�J����L��4'���J����KC�N��x�P��Uq�,z�X�*Q"���ȳ� �렟�z�+���~����#�����&��F&�?�5ߵ�����H���!���=�f�2~�k�G�a�(�e�c����,���׭Ii�����9��U$j�*Cc"��彂2��%��tv!0�ړ���%���Y��ɐ;���qK�vϠ����ly�x�8=���V��;��Ӌ���7�x��x�R�h��,��N
�w��yL����w��W��}�~�e��lZ�G�!������l�@�/��ؾ#A(B+3K�G�럚���8�'�zt9�oF��o3�m�� t3��b�~7zh�Z���դ���_p��si޻va(Y+E��ap��'�ŷd�P�̖�����A9�
���E�|ߔ��M���^�#&�Z�t@�1�e���������f�u|c(�ņ������M���}���C_�؈}]�}��eR;Jw�)����Nt��w=x��P3M������v��Z�)�4��Z�����x�f�<v�t�C(������벌��`��ò�C��i=����S�I��F7�M�% �>J+��@��4��Ϫ���Y$�gM�D��j���N��dq���fI%oD�Yǡ�s=�����Ĭ�١_Hn|��il��$��?���[A��,�M�������� ��UY0]'E���g2&�)P�kun�<0(�0 A �^��Jf�w�LTmE����
��H��x��q�Ix6b�f�!��k'(��!zЫ�W�\V�a�T4��֎�+Ϟ�(?�fL��T���>�CR����+��h��,O��K���9���������>D��z���j���sp6��daZBV��?�Y��%�V��̩S"�~��s�bsQH���;����9.��tx��6���(+�K���鹒����S�e��K�Ub(�wIa�9O�'pI�1/�Ė��C�Vw������4�= ���^~���5��;v>��)��h�j���G�?�Ұ���h�/vHźV	ܣ�O�߲c�m���oqR��I��<��S�GC๟��p����D��c�[az)�j)�"Z2��� ܄����W�/���k{�rM>�o�\X���K�-�t�YR�	j�����VL({EUt���b�<���E�4%ֆ��bk��t�S�@;w�P#�=h��Lt���ts�Fs�=�9�?̏)M]�8~�8T#�t�� j�>���L2:;R c�)Y=��p\��j-LW��j5F�C�X�v�3�PU�\̻�e-9:��m�$�M��%�D�zx{�&>�cf��[���i�Y�X�?�	U��,����[ĩ�H�ni�� ����u(�AOviȩX,�Ů�4{�$���Y =1[�3\�@�i��4Qk�@�h�;9+�[F�g�9A���\����/k�9c#@rJ�]���	ϑO�.�b��2�<��P,|u��9:�8������u�=�Xa��a,������=�ǥΎA�W��6T��]���I����|�r�6^R������FE}���D�XO��Ԙ���Lj��COo)��Z�D����0A�ݎ䜹e	�U��%L��m���Oi0��R���#�P�Y�>7�0G��� L����@��^�;~�/dr�c�9V�im�U'�L��ͯ������OF����r[�GK	����U�����T2�!R�|�i|�I� �,�p�+��b�~b�O���\�����5�a!�%�0wˌ�K�f.�����p�[�Wl��Њ�1�#"<s>��N�L��p37a�\}��&p�����І�=;��[�"�9��ײ��0
-�p�A$��n52 $cG1�#�$(�0WD��T�(E�D�cH���D��Wh%�]=����E_���y1����1��s�� ]�D����pևK�!��U����l�����dbHoeH�2�a�l8���k�,����n]�s_z���	�J�mr�e�zgVI��*�+l]��6��V����4�D�8��Y�)@�껜�b�\%h��jL#��gݠ���J/�&�����ʀ]��XCٷZՈ������8�>���xe-��NOv |v�t�7��}u����L��q#�Dpq�
q��њ�jN���T,Ǖ�-H=�]�xYSO�+AʹB}U���+e�ږrKF1QmL�Q[���=I�2�Li`�Bb6�b;^>�����&�7:.XHCf��)t8��vʁU�Y��4��P�B��x��/����n�c� ���b���]u��9����:��xF㇂J<!���/
w27b�`������T�����P�/�Z귺�f�r�������1vU�PG�/�K�������e�� XFgQ�
�XJ5}��K=���VS�rL�`����+Ϯ:h����dP��Vԅ���!�r�<��OZ�O)g�A	A0��~3yH:<a55^&�N��dĩ�`G�W	��u<f�Z��6�o��N
��/�@*�>:+H���B���O�~�^,[0������R*i1�vSW<B�;I��O� R$�A�+������oR4x��h��P�W��e�O7��^ق��_����5�3�%l��J77\��� Ko�+(��X�B�';F���7 F@jJ ���Ƞ��hȘL�3��?�r���0?AV�����Q˻�oh��W/��z�O�����j�w�fdȢV�_t�j�A�F!�۷K�C�Y`���wGYί7o�G�5Z��E#�	������!������5�m2&��B����A�#C��q�z��-���c�Sۭ#�U��*�(�ߜ;v���� �V�>�t�Ur1��h{"�?\��'��Z�Z�I�ag?V��;��+�j����:�u�$P���t�pN_n�/ ��J��'2�R,j��p�vh�����=�L~o�a��[_�Ec�ª4!���7劔1��+��*��@��?����uà/��?I���9g(����I���`�c����#g�x���B�����"]��� σnj"�:�Hf�Ӏ��>��lF-�b{��+����5J�<���*�.q�76�r��9�U;u`U+�k�tGٓ�k_d��M =���늗eJ��M�~�&s��Z��~\����63l��@R�i=���Lh�w���1"TQ��d�i4�:��i��s�W�ea���aq�0{��c݃hB�ૈm�����,l`�#�>Zԑ��ri����c�-�T�xh��X|�]Ӂ�Rv�]B>`4��%E�I#�Y��o�3�W�����%؃S �}<8�ϥTFЙ�i�c�����쏔!6c@*��ɫ/̗�`���'�`�jnE^>�OX��Ԯ�|��+�!յ����ߋ��;������&�z,�֓��9k��g��h뙚��7p}F�z��Lb�E���_�ꊣN��l"��+�f6S��U���.�ۑFAo��d�c
���;onc�;���gv�pP,�ɢ���34��)p$h�6�kO:�>�Π�����LBS�:KnN���V���@���%���,�@Ĥa��`  �MhX��K.�^�'m���J��(巷Q���W݆�7O=��� ��&~��db�<,D�Y� �e�֭p mC�I���
4,�\|�z I#�F�����]�	�RA%H���D��|/�=ٗJg��4^�YZ��T�R�G���e[6*�F<�?�g� �)$����ט�
^��i2���9�_ ��b�'F��0��:JT�1�F6���r)����͆e�gdH�����O���$�r������aGo��4?������c:C]�Dz����m�i��i���\��A�Ŏ������0k 
w�C��{=�F�.櫦#G�l�\�H�bXV�R<O�7� ���� vN���A�-:۰�Q�^�/��5_�%�*��fU�̖�Q@��_>��n�X��<A��B�����I:��*0h2|��Wv���@�/w�Nׁ"@:��$6�������+P[�B������$8�^�׵|mHC��%��,����}0���wU �@��]Tu�������*i���������6���?X�OK,�9<��:'�u�[����ʯ��:���M��H
�.��)a�{���T!��2$1&�,'v�l{\Q@̝�~j�@��z<5НS���C;��͞')2Qo��%"�o��b%#�+,�`z���Y��L2U������(x�p\�5�^���Z�ڀ4"�ɚ��d��4�ނ���Q3{8��!3ɽ���"��z>���ĄS�p)L{��]���}�"�?��[G�����%��Y�VNU�.~�"xQ���.��$�ydJ�Ӹ!��pey%dɜ1wpB��#&:K��෼s	bz��ٵ%�� \��x��w{!قw�YLE���[z��8���9�w�t��Se��/#8R^xr��M�iF��ɾ�ܐ;�t��l�4`�D蔆$f�O>��|��k2�����a6��L��8>c#�%t5ªJ�tK�'�=�6����L�&��p�y��(�xC��S���m�/�� �]2>���V`1V�l�����x� /��2��f����}�}�����͗�ଯ"�xv�NX�'^'��y�߾fԄ>�z:���t�ٷL���\Y�%g�]�}�;�|�=�]XՌm��jg��5k^�_���p�`�!UXY���5]bh?��OE��t�s�;}~^ir�MѴ��X��3��(_*�����-���O�����"�:*s��bDx�o�����.�y+�!������Z+'��S%k[*y�Q��@�(���$H{u��V�ƌ'���TT�PB�N���O�l�'/�t�<b��W�{��2n8ç@��ȵ��8�|<v���wk }�g�T\o�V��e�=�S�{ZSvGH+�?�f�g�xJ�m��j\���$������t�w��mz�^[[��@������n��<�L���m�(����H��[��	��
']�B�Y��g��J�X�,L�%+�H��p{{�1�Ӡ��zu�!��E��t����֐�l��-)U��P�q؏�C��)4Xm��wL5R�qZ��:"���mr���ߴZ��v�����?��u�� cۿǷ��D�[�-0���Ou�@�:ÿ�B^0 �^~N}�%ԥ��5so/RO5#������?�'�P��!�E�e�e�;�p=md�G�����^�Z�N��y�r?z����2��䏨�2��B�n��T�(�w=�yt���ex��uFz��i�l�r0����~��e=8T�I��I��?�O~�!9�eh�3�J�u��/�(�6޷�Wl�B��YT ��I&-MY���rrw�K��������qV�d�U�4ĕ!*�����1O����w�^fSӟ�@p��)1��4
F�=��eSM�!�b�>��Y�K�8 D#W�?�gߨe��e�:iZ|Y���5����x��+����CO�f�G/F٨���r��k��M�Č;҂T<���=�w��Zg4��!]i�0Jl��Z�K�q\�<���Gv���5�'0#o|�����Sz�ɠ�`�}x�C�{$;�s��f2�Ƣ�v�/	�L�m�a�p榁�/M����l8�>Ր{R׳�h��3����vn�d����g�3�1����	���H3�H9	���Է�IL�#GH�0tS{0`��@4h'�,��9�}��Q���wB�[�\c�nK��ny76�ڑCq���C�I}�!�Ε�8*1I���vr\H5�n��{���p������B-脕y8�=�6�GI�$<q�@?W�Ƹu$S
W��y�W�1Br�5K_���ft���@��9?�S�{r�M�ؼ�n�o����2�I�c?$��-x*�)�@�n��%�/^4��c�_sT,�..(=���zk,b]��Ձ(�іe�Y)���+@�#�+��6Y��UR���$�dy@/|�"���Í�X�%7���H����RK��j7=$���y�<��/L����H�z�@[���� �q]��ũ<t���~ZS�ce�O�V:��	_բ��au�H5���u��X�@��~O�*�2sͽv��
�{���Ț��k��*�,O�WT�4k/1#?ٮ����Q�n�*0*�)�r ��Be��"� ^�ɺu��mq�uI#X!X`�Q�k��'�o$rsI��ȯ#$��p��U����!\A�eًP; �e�i�FLm9���z2 3>�8p�[���i������%��A����+����'!4��UT�/ﻳ�w7�Y���%���#ݬ8�'��pM֪Q_�me�&�C��A��'*��-$>\��xj��9F�ۦ��ӡ�q5���:�p�Pڞ�+g��p�fe�����)cPl�� L*�c� M��[��M��I�ݍ��jx��!Y1k[f-{G"]�`�-���䴇� �����L�M8�F���S)���KIB�lA���.�d)]H��c���OVƁ���ݓî�%%!������	A��"��z��,����n�5�����"s�L˳4X�b�P��	F�w�Ң՞1-Z'��=TK`�.}�_��Ē/��{`E7_7�6�n���呖��"�;��U��7e8G�0��("¬h��D�1k����u��� ʏ�L7���+i_R��Z����YԲPV>ڇ�),�(]O�O�]x|�uĂ���D~h�a��
h�Ӳ��A>1�KC-��Жk�y�־���L���hd���H�~�ic.����;{�|</�A*#u�P��n=��̽���⮨i�Y��T/9���M���@� q��Ű���Y6��:AJxct��᪅��M�R�������0��i�{�~��[x4 ������oӜ����(�x�~�=m�[~�Ͷ��_F����l�_i-u�<?�H��� �Z����xn��a8� ��Wb+����KvZ�L�w����pA=�)*��bm���:�ۏ�e�l��cd��.�z��k=gz�*J(ݙT�4�9�U�� ⣄5<���4�A~���Iم/B�S�9������`N��6k���7`��!�������ۊ8�s�c6Ϝ�h�bB��i����W��d�`][����j]߹��)���9�� �=`�	^B�^v)"�3��My�Tv����5��z7@P�/rm��f���q�"�]*=g�����
�UҦ�����؍Y��f{!s�&v�
aj��;��wb.�"�#��'�ǧ�f!�B��f?[������!#�����NM�L\��Y�Y�AVG�Rz9��N�4M��>�[��KtD�0�}\�q4���M[`Qj��2�_�����4�1�I4��yk��i��vioa�E_S���w�*!U1�������~``�p�h���:_y� WI��^�ˀ�.��E����f�f����7�F��j�����nN���Ҙ(.��BFn��;�M�z`٣/��}�Fr��� bϔ����u��"g� )��,�^�)���CiF��kh�G��(v��V�+u�/&�:�+?+�q|��9����WGզbj�m#S
���iy5>�-��>ё��O${�#_����k��}�qT��Z)R�h^T�ak�R��G`u9�61���\7���#]�����c~�%D�4��/�')
�l�<�:�#%���V*m���u��h�'}�� ��U�lp3�3�bq4��G���A�35�l��}����V�w�E������7O�6�)�d*a���:s�_sFfЄE"h�ᚌ/�s�X���l&7������*0�\@O�'���e�{�,Y*$tNW�!w��������:�9s�n�^�	��1Dq����(	����]����S�6�wb����@'bcK�rԸc�*)�[PCkg�7�6����m�����[����ڕ�wJ�Vn �s�⛜�������'�`����q9}J��m���ߞU���x~�EQU�1�/dK­���q���wɀ��πئ&O�uf�1�48�����T���v�^����.-H���0��F39yq��m����Sl_�\��,aQ��KI��;�p�aDu�&�;z�($�*�����D���
�@.S�J�"����a;>�R9�
(O��,�J���'��!74j��a�HB���2K@R�@��{�ۓ>Q#^��i"A�wz�.��ߠ���N�P�XZ�1��ڼz܈)��*2R�l�=�0!����-����O|%T�ժ>��!	�(m�׵q�W�<`GZ=��_�k (�.�]�,�W���Y�+J�\��O��(0�y7�In�1��zֶ��Y�q���*>t��׌�!F�z|n�������Ԧ�[j�T	!���12B���oka�B��ۛ\ݎk���w�֛sL��p0���'<�ٴ�����(j�)M�فWp�H�̙,��!bG��O������=��55�˓Z&C�h���ͮ	A&�~��ɚk�w��1� )�.{��@��6�΄���dL@_��[�v\�!FiXAX��C�i�K��3Zh] .[�Zv8���	�F5���LS�l�	u�5)Q�kٛ�:�"z畊k��G��B����b���<ͦ+J�h�2���`�wn�17��x��q&qD�I^ �*��"����;�E��"��0T�J�8n�j��!F�\��'�Şp;cM�����|��e���vsy�UTQ���y�ǰ,�[��t�ۦ�]Q.�%�Sua	�������?�|�&Wi�*���@�|��E����[Ǟ;ȱPY.�&���>И���o�6����F=�vr�L�\)Vt��=ঘ�kn�K��5&��jZku��8�3��<��WC,�E�Y���vDׄ(ҋ$��=���jv/�@�c�f��Fuj=��k*�f_	V� ���'��Cm�p���� ���0;�܀��7�^�����,+��md}\���V'�h4-��tQ�����˦js����jn=r�1�m'%��c����7A�ߗ��?���v���U��n*I��2y��%���PC'#�F�?W��A1�[�p!�S��S�U)~�I��_�?�6�c��n	����L�!�|��\��1����+���t����h����?6����y>G̻%���Α.
O�M���wXDo���f�-K��N-�� s	�Z�Kʕe�w>�`�1ޣ�eM璯_�vy�	\�v��\1���׿����7
�<����N�y����?Z5�H !�IT-%g
�~�� �t�"
dQ̻�17?5*��@�n\� ��R� Y����@�m�dl��=v%�T�v����p^�jN��k�W:#I+J���`��.����k�6�p�X7�/w� T�Av���0'$M�%�ry �{D�Jq
�K:U��:��WN|�΋hO�<�`�����z�E��S�xR�w[%�+E�Ѥ���4���>��:p�5�E���
>a�ٴ�_�l6RY>��jF
ڸu�1�[`�c�����
*������� �v	�dK�9�V��H��y���hȧ��.II�X�D7��/%y�D%J�Sg���D{?S��mo�l*�g���	D��VOcg+�0������e��,�t��
�����&{����7.�0ݭ���6d�iQT��e��!èM��Uk)��Ϲ�_�0�TgBY�ʬ���T�O)t��NJl�h"��u�� �x��@�@"�=���%�%s���-r��>�1Qp�5�|�e`�k�w(�;�ׅBƂ�׆t���&+�_$�¦iUi��G&P�i��X��nr��N�N���Q��"��w��Ҭ~��p�jI2d��)���y�A��؜���9
O���,�aMo�S�ถ���%}L�Y�-��� a�_�e��:�[-�����K�qo &��.���Q��(D=��ᵙ�t��.�HG�_O�}�E[�CKA�M/�v�Sz��$GO�gf�/P�&l�����ni�X71l�?��yA���r��� G�E��Y���D�}��kN��U*I�8^̔+��ʷ.1�V]PU��V44{�2����I����`���FvdG2�L��F�,pU6o�wd�]v���І�!Ozj=с�c!Z�K��;� ���2�I|6�(�.���� ���,�^}*O�)?�ED��|��`��^9�L�%q㼙�L.fs��߁=��Q���(^�y�����9߄�������@﵁��E*c�ĳ�LE�W���$�\���	AM�w��FG�2�Z\%�;*E�֑cCf��W�T>�Fˉ���|RP��ʞ4��������B&�� .�N��1k��D��F$���-Hc⽈ˈV��"C��w2j������n��Ǻ$&~=vW�pf%�0/m�񎄊��b�e �-��՚X�+�����0�]��g+_T��\ջ0'�b�< A�mo֧T)�5�1Y���7N�N�{��phB$�5�S�zq9-�ʆ���ȵ���B韵�B֋�&O�%
)@�S���q�<Ff�����R��MA����UH[-����nX��:+�'{솉�rK[T��X�����:�'u�+d�Pp��p��1���2��������kA�B�͂ūn����1Q�g��Ʀ�e��;/��TZC��Mv������o���x��C��X<ܷ%�%��
�P|�H�?#���eg�+�B��g�ߖ2�76<:�x��SõJ������X�ēm�6��e�D:?����T� Y�pV���U�G�hh�E���:�Z�h���|C��V���c<JȪʵ£"�a��!�c�MGzU�o��o��� SL}{*�& �QD=vj��cb:t��MR���qE��H@���	W� �6���ciHɿ{�TjJf�e���&���jY��`���9̡���*}#����M�3N�UXZə��)��P\������!C���~yysB�J\ӱ�~�C#��P����Vywh��j�EgG�8�ǅQ�����^ϭ2g4&�|ν���C\Gtw{0�9���f$j�i�stk-h�d���,N�_N�:�;�P-a�]�F���P���c�B6{��6� ��4pa���P�d���3HĚ���(;3�H:/����5li�<}�����ʥ�]\�h�,�!t<��_vav�I-�(��U���:���'F��^&�E�}m��=2\�>\�����c� �]��_cC�l�CX`�.���N�g��i�p��^�b���Q~��
������	3�L�9��j���k����!�՟`����뚻ƛ���e��r�f�}q�傂-�����Z�M��D�? 궱n���a�!D���ɀ�����I�I�j���L�:�%V�o�AhE�|E��Ok+˜*f���(��j�b%1��q�q������M�pr{�4lJP���6��b�f�0��*5�� c6.=�=p�A4��:M�-~1�N/Wf��� ���8����3��-��p�#&v��A1�W��'����'
�������3�C��:~}���CaT<� ��x�
2��q��aAO�:%�mK���ޑ�]���J�4��f�j5�<pT���z��0���@��G='BY��	�u��F��&��T��uu�\<�����s���������(|�{di�Nu�o����'� ������'��׋̸�c�H�.*喹M��I�X�Vj����-��d@y�ߢ	��] ���xuGmZ٣�Ht�G7��/`}���Ĕ,w1Jbwި7�i����5��˦\K;.�$m��]�oJ���ܿ�S����M8���V�����:L�;��6�;�h/h��Ȅ<���GP	���x�Vׂ[n��j���N*�+,����,o�� Z�/p��m�����5�B	a�Q�3���В4T��CZ-��K2�(+!T�^��K���e70s��D�Pn`E��K7�v���7�eE�`�>��C�'{y��n	s��eǵj1�Y�S�,S��F;k���$ϣȪ��C����j��p�nR�b�H��$�'����'��%�VBD�*��@y+w�	ѯ(2�#�L�u�%X"����mi[���䗸�጗�����i�+o���� "?�83�Iya�I̓f=�/���X����sr���Pk�+*��[<A4(����Ŵ>��$g@ ���@�Ԩ\!|xӮ6��x,������v ��UM�2j�����jd�$�cx��iJ�*��ِ��,��x73�9�M�Mi�Ur%�=����U�;�D%C"ݾ�����m �p�ܤ���p��"�O���aW>g���%����L���bT&p���@kM�����uK4ʳ3�/���정f�s�-0�^��SDTV��|���2�<��m�l�_8@xe�߇��7�JВ7i���#]���)��[E�����#-e�wFGp�/��5�/P $���	<�ծ�o�]K�번y��e"�&��R|A`o��/j��{��x]�y�"��4HH�f.3�ɥ�u��)����G��O�6��1��&dĹ�q��4_X�M~�a�j�S�ooP@�hl/��kb%�V������;���n�O7�����q�i�4+%?~��8�8>�؍�I�bG��s�%�����X�|/Cz�$0��k���EO�������}�Eq�����e��#�ˍ�"�fv�D�@N��T
��ecN����HC���$�c#�?d��\3ho��ԗJ7�@5�E��+�ӡ�R��Qlg�j�[l4�h�
^ѹ2R(왔-M�~9i�1i��s�r��&с�V�j��ǥ L>��c2|�w�#��$��O�)��	�����X�����B WgL�~�����"��[ �@G;n��!R2FJ���.�������8T���$�R}����݀�=K�mXN���	59�hӪ�%8< zNq ���vQ|co�3� )���ҫ!�2�>K>�?-^!���%�w��+SŦ�f�CL�]��v�|b.���8f�R���XV��S�N������p������vq%�.bq�Ȝp��Y<����y�֧دԄ8��-L�a�ER� C�9����bޖ���Ҋ�K��k��WC��0�1���̿jT)&1����v����EJ�k��I�iCK!WcC~��*�� �d�OԕhrH����A
j{ɤ��HY���N�
����?�0���G�R	�P6f�gyv�ig���BVIB@���+���Fq0960���k�B�=+_��i�u�g藪%�2�0ä%_%�����E){�Gf"��R�x���S�I�풦�ݍD.o����:"�b�@��W��>��X���|�^{)_*��FU1�,'<�����i�8�)�*Q0Q9���=K繕q�*x6V��з2�:�;C�xq.�J.��S