��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su˸Y��'��d�Ay~�`�i���o3 1&����1\T�����	��!mF��
��\�ݘ�#X4|'�~a	N�1�""rϗ��?���ݝ��^��lt����d�k>O@�0�#/���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
N�m�H2
��j�Y�?	l�Aō4�8�����>|�f[؁���
Ζ{�����0>��������'l�d�b�%#T���QOo�Rh��&42`�-�R3Ml]�Gq�]O��ל��J���('���Q�5�.����p��� 6�	J�/FM��8���b�)f�ĐI];�^�EL���j�����D�1�5�1�K%M6P�]���*"&	а��u��~ٷn$5h����k��O��L���׎D�y6"�  UD㍺���"O��ܣ2^ �4"�.��d_y&����V���k���ƭo����`���%ȯ��e��εA;�3Yй3V��l%U}��N��������aUiJ��������X(7:�_0�Ah9�[��=�2�5�����,�_���i+���C�m���K-?�qi�b<�-�a�!?@�3��w"�[^�J�������+��A��W�P���
�sYy�ŏ7j�S�����h����nK�L����E��#��-�\�9Ú��U���-|{s֒Ѩ�y0z�]�C �_@Jn b�K� ��A��a/�F�B�!�Ma��Y'�����G������]�LQ���|��gE���,\6���Պ�E?��d��򄻙���R88���Z�c��5���G��{,]n�M��������ܵ�l�{h�W�2;��+p�εn���>"q��N�G�T�����o�-�m�%�xG
�o�]n���	l��'��a��qB�d\|���Yc�Z�t�x�塳Lr��X��/'>]��59֥�'�w�ƣ����2I~ٺ}���Mw�q�ckg�<�B��<�� �b��ű�G̹�[�(�R����Dz��#hu ;��9�`6.z\��".����X*Q�dP�So�4�K��z�~�n�^�a��W��3	# ����k%��t��S0��9����N� �o�����.�Nj�z쵱�G8b�1?�v~�W��e�POOs!iъPU1��� ݀���e7��o��^�]F=c�59�s�+7�ҫv�J7=���z
��_�σ��y�\���h�_��s|��Z.����*ô�XE�@�L��:���e�P��E�U��2���Ἒj��iu�*�9*���^�y�Y��ja�3����qL%Q~����P�l8���Y����3p�V_�X��U��2�p�R�
J��p�ӥ�-�؞7�;���
����ԃC�B`)��Ђ��#�L.��FbOx�4��w�6�c��Y���ia�W�le�\�L����
NBR��@9��+����dϜBF�5��q�>��&�.{a��n��k��/|�i?ڜ��J���|�pP36���ҕޥ+�ϻC=�;7_!�g}u_�]�(��1Y׵��B��r����Z���aqB�������_��2����<�g�$��mִ�Ga��)�f�"��{(�3w>�R�5��D���t��8���A�����VkQl�"3����}�� ������z�����T�Q��@f,�V	�
�ib3-m�''�)5�4D���{�c�+&'��'�}9�5P�g8�����-;iaJl�$��W� Cǳo��zH��%N=����Iq�>n�0��| �H0�,�X�RhKM�Xۇ��tQl����Ge��j*��x�G��K.�"�b��.�o�\�����Kg+T�Z�����m�Ĺɤ�
��ó��&��)5�&�+�m,5TPY�Vw�~%8A|��=�H`(���JآD�ދ�(�K{B��ҝC:�%X�?� #�4K�������lTH�C˴�t�ԕ�(�<tۋ�$�� �?�R�o������|����O܏0qt������4����/a�+&[.b&����	�Vo�-�0�,�ɽU��-A&4�#[��u�d������y�e*��]�E�����1rGz�D�b���������?��C`�� �̲�	�Į�j�>|e@�T9�K�q-�C���7���C�kcn��DqZ����!d��su&���������}�[����Y��[�m��%:M邮>�6�F9��Q[���G�������;cX��S�/�n�ug�����y.��ዕkkc��=�w�cqsܲ�� �ڌJ\�_�:��"�����w�Վ���������2c&S;����t��v��<�8��P���hhk��,���%�z ��M6�a�s��Rp��7��cѮ0���?�Py���Ada�Q��
��:�2?��B�_U�Q&�-^�&�P��u�r�hD���K��8��^�O���O�&3YC�3
g��S:���|�P	��E8x�	]Ӂ�,�h�����s�=�`<���B�����x���.Q��l�5��U��t4.U�`�a� ������G�񽏞}��qN���a����YQ�Jl��&ủz�$x�X4��3:�Ҹ �Na^ܵԈ�<ME����Ӓ�P�k���~�[���V� �J�i����z��`D���3aתH_u1S��.�
A���{��(��H;��W����2��W$�����(���6�ǷZ<>�a{�bh��=/�	���V��"R'�>�n��x�Ērw��Ĵ\cw��]0�Ե���b�Ԧ%�8�q�7&�`��XG�ʎrqL�^j��O<˷�0���fU�
�Bx�,���b�q�ade��h6�
�o���O�����{U0��)"��ɍR�|����O��4(
hqµ&�]b���T
��i? >+'d��GWt"8�I��8��8=�,C}��
���G��xw#wj�2��P眂&v��aEt����ͪqxJ�� ��`!֍�DĘ��.�oU�F�����m�V>ݲ@��%⫰iX�2�ȅb����-* �0��
�%���P���3j��7���r ��<���-���_>^�����s�fs!���������;\���:�R{�f����L�@�c@��p���K�3U����*������N�/�p�e݆ư���4�c.{	����yJ����4�4���$_�>;�ƖɟQ|�ܽ�zVŬ�a�����"r$'s]*�.�o+F�����*�\��8*��"�+�M@/�d�ڔ>/���])X��������7v*�
;�
����N'f�@Z���k\s��eFz�'��G!�>Y٧�B���n�u��Ze�I+�W2e+����vhr��kz�S�[�E�I��'�1����1	0?�������+�GhZ�r83aA7K���"A�J8��1� �t��L4�/��	�߈�",Sk��t%D[��aF�u���6$��,��d�D]��� �J��39%��J��`z�3�;0���|k�U\b�a���^�M�:�ݪGi��_�6:G ��y� c���e��R����.'0k�]fw���'If�aug巀c|�ݩ<�dx%�jK����<��t4��0���/P�3��%Ѭ�;����]ʹ�Z��I_��P9 
|���,�9]�� E�t��($�'�gE^*X`�\ v�S8(-\� �q��5fB�w[�=u$�.i���Pվ/��dye��vDP��j%�>dr�#v�������ׇ��o�/��b��ʻ� N'&���H��P� �5��Ot�q����w?�D��_k6[l[�8���k��3`HE�,m��i�0�./�%2_����P���M�����P|D�I�J8e�� ��e��u��Q�h��3?��vM�V��	�7�����q��;3]���U�bC��Ѩ��Ps��3+��>�Z?���#��PE���ǭ�à�d��]�PbD��u�cC)�iv{��>G0��"���+]����'b�5�����w���B Z��i2��W�C��7��:� Ȉ@it}�&0:L�	G��c�.'��$>��k�r�8�s�cT���~x��/�e��z��ז(8�V�ǔ� ��	D%t]�% F�wt��h�JzY�(}J{��lW��U�.��,e�����$h�bF��z�����OP�y\�p��Xz��tj��<�[�� �H��X���W�#�#˔�O�-��J�а�ֱ�� ��}!�L��R!b�0h�r@�^�x�1�3Ļ���9V�A��;)/����z�֐�qTAnF>�1�Z���8U� _
��!C�v����\%�]e'!H��%��RFV}�s>��*�J4�_� �����*aXZ��$�QV�x��gKk5=}�WX�ԉcz��U@�"lf$;����8�A��gc7i"��<�16�����%���\�]����8q��S�[�Q�_5)nۦ�V[��M��4�=��P������1ů�>���۠��|Y�dv*����p'�-��N�X��nC}P��e���Z>�*��K�=)h`���f�K�������5u���g��/RM����G0�*��9��[�~7G4C7�6��x,�k�T5�s8� /-�>&~��Yv��П(�>,Uo@6OXd�0̂E^�����⨐0�KLX#Q� �P�m�8�ذ_w/�,�3?kȅ�Wݗ>&�Ǉ�7B��Pl��������
�IHSFpS��W�m̱��n� �"�QX�lJ��]�����{���4�g	�`5�-����a�>�nދ/G}�	`cMR��Nu0%��v�\I�ê[�#��&
�}tBt���0�6#8���E�Pɘɛ��ԹS>MEi��W���lXH�6�X�!�"���-:��y$��_�sQGT|�+pȾ	�ɀ�XK"r���t�����d�Q�otIٴ�Nh���$��ō�e y�B�ᛊe�/D�!�	~yB5O\8W_4O���p���;��_e�0;���0N@�k=���A��� ��I�?�D�O���ۀ�HR�����2�N0���c�B�}b��?i̼d,=S:�!B��G����q;�G#j	�S�n��K�K�Ծw-����Z�����@�E (�B0�������U�����d��[B'O�t��jx�7����b��~��i�% )I���I`ǍP7�*0K�?��chJۂa���Erzϕ� ����ƥi�25x�e�%O&���������6:�=����bE���e6�������(0��Q������Q�	閆���scZhR�Z�a���X��]��\5�;�Dw��{
�H�9��0�%�����>�u�7���,�47"�+�ɇ�P�b͐���}|7v�(���0AV�fΚ�O�������7�Աot��Y=f�4�N"�����֟�c��yQ��t�E���/���vp�: &�ϻ�����7c�F\��KI]��S�p����`2�^fls�E��2�=|�U�m�\���ES�����SpB�[��^v�k��Q���F��׿�/x���W�v�򫧿ǎ1�O�>Y$�;�i�ܤ[���>C �#C��\��"�=q�퀎�iE�m�Σ��]�+Xd�Tz�˧n;�TѕK�����1|�8�dZ�vr����FR����h���G���|C�VkP0K��F�;dۜ5ߙ��-���&��D�C[�sN}x�.b����J+�O�]�������"L4�͖��-���KX�q\�9�����& �g��*|`J��V����'�i{��{
�w> e�Vk��|qG�O��^����D�2�� �_�m����tBg�UP$�����~;re���oH5���I�%��}���G�h]��W�i�crsO����, ��9�f���!%^�%���0!�S�\���m�;pS[�P(8 	jc�T���A�K��	`/�ۙ!�Ew(��F|B��J2$��T<�)����?,���U����)mb���l`~��W�S�gA�Mc��
��g��n�ϛ �"3��S �y���(�@t*��u�0$���@�Вc�����L���X�H�!hm�F8d�
#�:��w��WO�ďȄ؛F95H�G�l�׌s��\V��w`n�\=�auI��<�Mq_��:��S�,2�7R'�ئ�����A<�IqX�cɵ,vF5�[�sB[A#��������}Hj�����WZ�ʬ���<�[�R��p��?�cgx��Z�Mb��?�����N�^���Һ�iC��I��h�̞�&��_}��*��Д���E����GS>1�������i�g�h���~~b*Sa�\Vyqo\�}�Ȫ_<x@�r6�X�ٜ�Q0(7.ƛ�����<�0�듼R��̔.�=�R��n�qb9�\0|�OOHS�^rʤ��F�0��C��z1���˙�4�D��gM4�?��{��s���0��xu���VN��y}����KUN���D��[ʜ��|�pLk�S
r��g?lH�/���%���梅,�kt�TU����7�>w�����F��o�G�9��:%�H<�\��1������?�*:����j�PL̺�o�����B�uzG07j�O�o���_��S�u��:
R����zn�a���K���Sŀ��b�T�� ��z4;���t۴S~��͔�$�����}��M���Xs9�bP���������kT*I��!�d7ؐ�����@���-�Eߣ53��yc^�����I&��,��дˮn�YqAn[����l���K�#��2�9	.��+(�&�F�P�j���Ȗ����H�_�u�=�{��>r0�M�U3�ֵ g��:B����2�em4��[K�S����i�5��s�ģ�X� �Dw�?�l'�f���HApqnӍ:j�8�s�Z>*���[�@O1�����~���iV�3��.�uL��U��@��ФSPA��v ����
������n[�]`���Λ�����4�ȭ!�F��;�T�`c��'��+�f��@�Gp��ۀ��CB���?z�H`/�
���.��˙�d����0_�M/ ���T+����0�k��oh�On޼6��a���Y8w$�F�����tx=��]��.��̍-x=���LU���5�h��]�@�ڴJ2f�ȥ�HN;�:5�
|}ٕQ@�C2�NL��F|�De������`��Z�'x�׍[/�qM97c K̲��e��&3���U����oe"��&���P*L������ �j�'b
���XFIsK����|���J�]wzY:F�z�G'�gc����Y�����T$�Cs������ʩuri\ط]v���<P���[4�"\zEzƦ��^�@>���|��/R�u,E5S�A�������X�W+e�
0`g�׈(x*]o���U��<��B��O]LaP׽��M˷�Gh��4�!.��	(�Y�ut*�I���C�W>��i>��,�#C%�VZX�1�ꂀ"G5s�@r&��B�2`��n�� �YTYBCf_)h�d�	^�v��ĵ�Vy$�,ԲRPj�B�/��Xc�o��5�R�ub���\�!�P����Qi�i�����ǚ�l	�b����THqѱ+6�����"h���pe�g<�BšA��`����	��Q�Ҥ����?�e޾�m�6�M[��$�ݮ�G1cPxQ��J�R�Tk�Jj0]31
�s@�;t&;r�E�[4·��WA�[9{pqӛ��箰�A_�L����\�o����vﮤ
/��'!�m�8�"�+t�!E��p����Y�[�&��5�\;A�/����eKr/����L�b\�ȵqL���u=���76����j�����q�� ��֍�%����H������� �7}�� Q��8�%���v�Z�/�����G-�9��U;(�i����
���GO�%Կ�����$��˭3^k�g���� ��Ԁ�"��B歫�!��U�u��wc'H=:_�x��x ��u�g��9���[�FY��Q�}�Z��L_��8i]�PrxZ-f�by4���A���2�7z�җ%�9�cN��b�:����Ð��\vmk�ؼ��m��T���|��ꓩ C|ͫ�>��.8��������h������!=��ڮbQ�]Ceu�"��� 1&\I%�
j���k2l���&�����x�r)��b� _�ΝEV��X/�9nQ�#jD���aŠL���>�jp\��S�����aB|3�
�{uй�YWM#�K/���)H0Ol6�	./!B����-�3�-�VϽ���.=�����J��8b�
�ѧ��꿞v%r��Uhd֢X��^�ˈr��z��сF"Ȃ��N���s�Zf �Z�Q���u'���h���#�6��J?j�Ĵ�<&ʭ�[�G+����>m�S8���]yp�Wf�<aY�ͤ���91��҇��vN+�E'&k�k]���s���>�S����Iv/D6HƀS
�!R��ϗ/f��;�-�Тꢴ0� bd�T�_�xz��QuzEt�:�O���X˄��m���H���������a��N�ns�P���U{���Υn�����@�Y]�~�7)�qW�(�p� ����E.^�ݼ$��:R�7r�(܋��ú�������z�:�tj�e4�:aIe|���e��Y~ �V�;�.&��(>��Dc���z�M$w{�+�3��_3�����b#{.�.<���#}�e�����z�aK[V�-c�E�֋��n��U]##6,p6T�x��ã��C�,�1c��l:�"�'��Y��Kت{���e��� �x�۝�[��%�vGl/ ?"�;�>�U�St�T��Was�A�^#�o�.?�I,��(^�dLq�f|KZG�;�a�Ӱ�7y�u���
�U�0I�I[�Y�L��^���m��&\$��A�(��*E�[�Oݳ�����e^m�,�<�[�:��cԡA��Ϧ�7�,�8�>�"<;C��6c�v4	�k[",������������t�Ř_����:�ѐ�~��^���Q.���TG���F8k9C�ƛ�\"���z:iT��ՆD���,<��o.�"�7�NO2���d��	2�P���/U���V�yrY2�;;�9s�т���
g�1/4G�"�t���~I���h4�cu�����{�����S�@0<ګ��{<���P�R�4���^�%8��R.�V����sboj�аl3�q����������IE@(��,���[v2�'��`����柔DEǯ2��f�{d�>��,"~}yd�{�:쎲�H7P��b��s����I�3
8C�?u�(7���.\���NL�{%��Ra�M�������&��Ô�g!�!�L��b@B���f(�����(h{��n�}z@�!���0���[�S��
�g����y^[n����(�d��SO�ϛ��$_^�Q���\�&�P�T���<GRL��{�:v��2�2��� T2I�w�&��~�?-qw�GN�? ��"���d)n!ܚ����X.��ŀ���J�:���ǾPk��
4m`�=�A�DX��c]��\Gӓ��3����l٭a�j����gz4�E��r�)!-��W֍c�5M� T���"���3��QD��0Ѯ���-�x��Ӵm�q�#��Gr1V$�vL�E���V�B��]�4eJM�ɗ"*�y���e���_�xu�|a���V�.�`1nE�+\e"������+9=BR�~�R���`��W|�{��&Ԯ�B�;p{���t���4B���h�[F�+O�c~�"dѪ܀~�L��R���b���j8?Rq���_�)���~�h�F$bR.U�ꪷx(w�d���Jm������
�P�e-�<{)���R�f�4zσ9T�g탣�A��8��_�w����Ӧ�c���wf�C�!:r�^�\����Z�?"����i1�]�ලP?d>�����;G��Xɋ���ϙ�-�(�n.�P�_X���U"��I0�dy�BO4�oLF��јփ8$�ݲ������u
�idH�qvQ\�����w��W�2��\D2��Z�Lx��AF��̈́�zK����� i��QHFUG��=*�[�M`ʐ{�2�r�X�~���\�x|�y7Sf;�<O��L ������Ge@,�Y#h��%�%��#�;�b ��c̋�<��@�z1Yb,��40$�b&e	4԰�[kq��0tp=��	����>�U8Y�G�^���
!=�^�ڃ�2RKo��)!���ǴG[<��1Ti���xZ�?�bw?,eA��t^\>�F�ƸQ��U<��-`#���]i6u�s8�b�ye�z��إ����Q�y%��6R����T���'�T���q���-�Q��OR�߸yq��7:?M�����%]I��L�',?�w,���F��}I0��A7Ŋ�Kkp�P �CrۈK
�����d�8T�|���b՘�R�w:�<��e<!>@p����+���|I$�>�T&�fz�F�F��G5���X"Bv�E[���r��*6Ϙ$���GB��~�wo"��'��`�I>K<���l���\�� �r���h� �ZQ����v]�^�ֆ
���*�[����o���®I.��9�b�c�7_�X_��qW���~u�Ax�FY%�;k��o���37�4Y("��1,��������&�w@YB�"���o�(�9�.eq��	"Um�ь� b|3K�恨V�aFܢ�!,ħ3�I���;PĀ���e����"�w�&��:����ƷO�_B��e�V�n�N��x{1뮗�1<*�+K�q��-�#�sT�"��{@s���dw��Ԏ^��'	��oAW
A?[�B�g�C�'��m(�z� ��w�+�AO/(��N�,�e?��=����kՐ��-�Yg<+"W�c�>�#��_
�	��<H��3��M��R���	ԁ�&Xs��:�;����H�Z�]�H�&��ť[c%�Z4~jӿ<2������ߵ���g#ǡqgy
�E��w,�D��W�$p��Sd�g�y�0�ZO����%8�Ql4"χnHA��G%1NvG����I$����~ I�<�;�{w���=���a���CNȯ�^����]�Q�=�l' 6�qo�C���Q^H���Ǩ��kӛ���_ROkݶpPP�}A���1[��l���H��.&q�,��,��E��b�B1�8�B�҆���Ne�1h���*N�V�f�<J[�<Q0w��8-���<�5������$��;�|cG��O���y$pe��"M�Qդ˓�IN�.����Ô18R����t���N�4�d�j^��m��?��I�O�����*[ ����9н�9z�R�d��%Q5�q���8_ER����d�O�M����n��0@���U)S8�����m�mDhz�?SJW̮g�D?�hu������ ;�~���j�A�'>��r��O؟	���N��B|�ۘ^Q�P
b��C3�R'z�.1�D9K X�U �u����J�N���)���(�`�U&�� �z��K8�	�~=,�[r�\���S�c�ߣ�td�dUu���n�.��V ��^!�2�e�r�.�P��dEU�ԏ�{�����S���p����s�������q�+�v>�4������Q��~�ѩd�nĀOOv�Ru�����/�j�\��NJ�g�*=��=��%'݉za��,O�g����@���I��-i�Z\J�ԙ
�e~�Fq�D��u9����+bOh?�)n��|%�lJ\��D��}��C
=;y)nڄb��@F.��e��;v�B��{�sO�E�;�^v����P���Ru���҉48�_@�
�H���Ke*u ���?U��Մ+ �2q���U�FO�����ġŶ�3����]��XDv���b~�߅Q�Űh2��2��ʤ�`�p�J��M۟�n�% �:9�{#VW�_����kM��в���4^�����G!��/���T��}��[3&�5�.~������n[7Ϻ��P<��٣�Z	���'�ˉ�o��F�L�k�f���1b�h��Y��ku��bמ�y�韛Ew0ZQ~�Ƃ��*�3O%�`H?|����q�&�]'�H.!��ՕϘz�`�Z�n�cpX6��޷#�����`�E�"�����5.s���;�~Q�Z偢W�M��G�W�\r`��)�3�}���wql`Az�)����{����}��Eg�*vW�W�pI���f�������c�烿��^�<+���R����b{�q^<��$��md���������s�������xF�ʓ����fA����;�JL��jӝL�� ���f^�[�r��1=b����7�-Ꭴ�$\��ȩ�N�5?�s6�[M��Ȼ�58>�������-��+�t>Ǣ��E��Y�A�Op���ނݾ�@�f�9�d3qE��s�oYX��#��$��*U���p禅�4���sS�ҨxEO���#3%�>����z��$���C擠M���(�C�v�Hʲ=�-¨�/Z*��&����t��jN-�A,J�9�(�]E�J|�6J�+�����wK}r����dR�h	'�H���%�����g1�2�+` Nl*�r)}[N�7	�xD���I�|�Ԯ#�aU��O�i��������	�dE�=��B=$���|$�:�^�b�d�i<��b�h����-J�@�.Cnqn���J��<��'�MC;������d�5y��!f��_	�e�G�nE�Z�Ao�z�j��8���&�R;��*���^���n*[F)
�c|T=d�t���aow��\��Q��'�*�b�C�xi��)�C�ޠ7�~{ Vu7l6 c��=��32ΓR�؏��}�e!���Q�����_����,9;;�EH(n�cG�#�� ��7o:@5�I�x["(NJ�:<�aL련����E~~3� x��B��s�&��
a�P}/V�qTɺ��[��or6���ֻT�~+�� �	��~�trڶL��~X6�Ȇn5'�D͖&?y�C�<�+�^`�/(Ja�<C���y,�u;*L��8MfN���<�KJ�z�_�����n���kL�E�Xy����$;�b3�!6��b�KDK(�u��v���>G�e3��C�묥�e%�����<�7�4fB��S�����3yIۓn��ji���.8]2�͸ۚ��N���<�o�ˁ�匟��Z�q�׮�b��o�.Xԏb��yԈ��,��_~#J��6�����L���x�i�y�f��k	@��MG�������)vSƆ�V�Pb)ވ �զ�~�~�:X�pf�#�1T�w(3��ǿ�{oF��Dd�-氉g=�\�
c����<��#Z��3y��]{I��H����
�Ko��W�"b�WrE��m�|>�͆�M�*�[�S���I�*�+��y!�֧�v�ς���*y�aE�>k��o��_���?䂽�>��	�K�$�\0hE�Zk�tv��7���3��9�(����!ҡ���6}=O�5�h����|��>��/q�nr��=�oc���c&v+Q��\�]{9�(�����,w�賌�a���*`B�C&�˖����sz{���@|B���&���vS<��ǹ��8�^�Y�d�ox��\�~�.���!#>$���Z}l�f*Oُ�h�^������f�����0�I�#9���'Vj�a�>N��j�6\`����P���6�m�VӿK�L�����o((�~�su��#߃\�_���~�T���3H���q��	��{ƾ��
j�?�vv>�F�j�9�?�.�m7�(����kݚ��pfY�Lna����G��g�R��h�����F��VW`w̷�j� �|��ZSַ����Z�~� y�u�F��L���@�x��X�� .~ZB��o��
g�Q)��TU��Bw#1|�y$TD��P��J ,r�ҽ���
�DQ޳�9��j�N,��
VH�!V����7ڊ�;�����R��\[�����y�|D~��m��7�x��od�q:
��x�{Ӵ���!�T�Oj���c��vq%i��⺇ٸ���@L$�&��yt�@��)vL���.CDXP=f��:��t��(�\,�"�D��q���I<دWz�x�������}�v"�j��b����cr����E�j�WS���9l�;Rʆ~ �?J$�%e��{._2>Q��s�mYc��6�B��v�H���q���:���X/0�!��pH��:��t�7_��aP�T����8�+D�q̈C5i��t��w���e	rۻ�z#�&r��x�E�e,�yZ�n��(*���8�G�}7��	���!i���n#׼�d�f�w��J�i������9Z�\���A�+D�\h�,e㚾��m�5`Z1��98����#�ߞi��}�q���QY�q��p��At/�a�XE ��,��֬��pkR��y`��X��kt��D@*
k��|��A�Y�+�Ԥ0�v�y�?�Xz.L�e���`}Jr�|	`Or_L�1|��4D��[� ����8������s�M��}]"���v��P�Z҈�	Yעo=N�ѣ��	UF�-���
I�WF��M�����D��qB=s�ǵ5�:���;V�Apx�3�T�On�1kJkN�>�I3G7���F�D_�e�N^2&��O"���		�/I&�|Ѫ��l��^w�/���	V���~�������ʯV�6hV���0\>�g�Er ��»�]��u}(=�x�+����8���\8�G{�B튆�N�.k`�l��t�NT�d�G*�PY�������N���X�*Z����9�6i���9 ��'�7�v����br�KI�@Ϋ�?�}5�o���aH��"�<1��4�*;n���ҙ�ۘ۞mL �އ6fa%4�0�+��y�)I���?�a���{)q��q����@I�	W�P�	bx�/�T��VfR^�z��K�~3�}�@
�>R������t~`&R��/xJ�X�eC�m�{QV])�����cX�HN�������[9��[�-���\W��c�Ko���a���"����SglҐ8 �D2�*k�(B�8��*������?�����@�Y��,|{4ǧ�zB���^v���+�]�g�h�e�e�6��$��f���N�y�Vn���}�ewԹV;'5��vn<z'�{s�;�����Z��i�������Z����J�_u��f2F9J���R\L��>Lg]n�N4�3IB��L"v���>#wu�b6���
W#a���P6���w��;�݇sڶ��1;�Xy�µ	�E��3�@}�Ņ��*�*��\�6��C6HO�w	�EN�9�f�|vO�0,����YՒg�>k�������'i-,�.��P��O�������[�'S�@d���V�ӝ>��DDTf�P�Iy0��'޷�[��;%N�T��.��_dvΙAJj�ʙ��gh�@,��e�2��^.�]�^1�
�ޱƷ�;�;8����d���'Ps�Nc#�\n	����\��>������P橴/�\�Kx�����@W3df���V� �|�6�S�nAj�G���}�.Am��ROׇ�ݬ���B�-�����!�L��S���5��I�۵�.k����)�*I �	��Q�p̵�p��ٓ}��������?�v۲x���F��ZL&Dunn��N�veNh�S6L��զz����Rf�wi��h]����s4�AR,˜����B�>�M�4Z�	4Yrl�g�ID�z��/�޶~���r3AhZ�z}����C�f��3#��G_��#�/�D]}*�|G�
e��h`��_��bl��nm��8	��7���7�)�V�5���]*7���<�T	E-����ő��\u�%�!K�ߵd{"�kU�dh�O�{āo/g�[��@�fv��P:�*��lթ���Vjㇳ�J)N&��y�5���U��Cߝ�jfٹ�U�����rj��Ҋ�~��:b�6ϸ��tnR$����T�~�U,p��I�d��-+����z���_����=�Y��;��� ���l��i�>���-2z�7����f��V��5�"�"��s�CS��� q>�V��?ԋB�+�0K��1�R��c�����ri�?
ߡ�m92J>gĞ��b����[��a`�Nbz�<��V,�ffr�>��˪!��0��q�+^�py ��K�n;i��}��NS#�!a+O��
��dV�QSFk���!W*�H�BH�'�Kf�p�x���b:�#e���"�٫�R�Jd0s~dS�?��3����x(d�t.���}�c 4�O@�,�%�������ISپwX>j�S��WKjG1=0���+�&���Do-.{�����Q��,4~��*<G���H�X@�wN�����a�� �uw���01��1����E�b��Mz�'GO�|���t3yG3d���<���XN�1ȰŐ���X��a����k8F���[1�n��]���c)���O��[�������$YvӃB�I' 1��Cǀ�D��x� �Ax��[x�V;��"P>�5��>s�	"��ٔ�Q�FIB���/��a�7xF����W��?A��N�X�$V�˩!��v;#�W��*�AIq�,.kdyv�A���grb��ʲ���E��9-	�SU��������r�5���FuT|��'f
ƻ�������1��`�߬��Qw2�D�}֮�Ot��n;���i��WC,U�U�;��J[pN%�R�}��֦�zCB[]E�B�c��֛��!��,[�$��A����fO~�y���y��Rl�F���Ȧ��-nOhB�n��0���c]�|}vn)�O|�E���w�(A�n�R���,��x�I
����f�l$I�y���&5A[����"r0pv9;r���!��E�l�{�ӻ�}dT�Zj9DbЏR��p�����>� T@V(础&mN�������{qk�(rG�eυ^Co�K���=��{����"�F�f��J�����I$K=�����͕;�g���&a�׿�B���Ƴ��l_�׌���\�S�ܚQ�VO� ̳���;��1!;����ZT��X�8���#>3U>�G�r��������3����K$_?�{�-H���NP�"�f5VL��o��-/�����*��!�r+Q^sM�S�u��uN��,v�?ٵ��ug�D�U���ь�CS���<d�3z~2�f"����,8-����	w-�d�vQ p����9�v�H�+�D���*��
�+�?�waU� ��ڐ��%@%�f�p=�0x}��&҄K��Z����V�}���$� K��܉R���ۆSHR6=�k��QS[ȩ�k��Q{�,a�oc��[*�Hz��_޵6�.?���t�t��I�t�.qm̬ ��h��t�un���X����QG�p��b;��%C�e�U��=[�L��Ջh�-�7L̚�S��c�f���2q+��Vآ�*�
V��|�F�bc�ʂL;�
���w�0!�0�?Ŷ��d���HLgt�Ju"�n���d:� �Z�\�c��-��O?�q621f��3B"�ȧ���&�&�����~�{�(a���·A���٬1P��6^����,�sK�&w�>Ɓ#P���yW�`{�m��{�