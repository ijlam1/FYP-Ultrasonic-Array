��/  �>"s��E��b+��	��zKœ5W3?�f���ڽ�u�7t�XER��r�����r�e�F�#��FkI:D~Zx[�ކ7½O{u��/V�oM�{?���lI�?���Gy�,�eN|�[:�ҿ��&s�cH�6�z���5S� ��r�����#��T�7	3i�;���FpoN�9m�̵p4�F�6Sֽlq���cf}�T
�%�y��,�f��X+o�R�݈ټ5rX�I|�i�ª���7��f'�0L����]N�Ȣ�3�f(��d��W������JA`��a��_�;n[����xЋ�V#�"�;Q�����~�{ZR0�5�(��E�TR�`o�Wy	r|�}߅ls���W��y�N���;n����V�k��=G��q{<l-8��3�B�>ǏyP_y(�ڦ�|�z�s�EK��(2�b0����@�����WG�>�iv ��v�?W����[� ���#w�iO�	$~����T����G�w+!���sج�b��O�:����L�-5�������]�p[��{�#��	���/u���M�#���eὐf�i�X������ٕ�v�i"]���@�a�۹�B�&1�)	[j1��r�,�n��[�V^`�A��֒�b�+9(��ohr���\��_�j�'Dg<2�my��5\��?����n�VTx䝅6ժ,��@؏||�F��2G�"�W7!��!.|t��h��aF�o쀌�B8�{��9�܈-�m�5�Z�����(i�Rz_�! �e�R�C��_B���f����X��7!��rs5�K��^(sJ��]+��ف��.#>����Լ��S�T�2�B�4r��kH�L�����������3ovٿ𲕬~#��.�����m?����ua��P[��d��>�N��O��b�T \��ḹqr�'�������4;>ͩ҂���e.�]���.{-��P��B-�{@�"n�K���}[��z%G=޶]�D�!�S~)��KΈϣ�Z�h�;�]>��j`�7��O?�j��B�.Ny@ͧ�����?�����tD�Y�d�����}�Z�U��Y��T�8�~R�~��p&�kf���1�Yn��N�b��;�����9C�w��̋O�t��ְ<k�*2�,�U�&$<#���[�H�iB}GP~ZV�'��ydT��A��` BWg���EO��u���b�x��h]�A`zC|R�}���ѲT�qVxS��Q���i�+�p$�Mx[5���������d!�Qj������q}>F��&Cn�۽`�X�+�˧�d��Y49t&�b��"z��I�2k3���,,��[O�\��G]%��'�ImG�*v���<��^Oi��f
{1��FN�)@�=ʉ����^2f�	1��Ed<j��ԙ�
Kh;�%-�,O��|��Z`��L�P���xr?���	�T�P}�R�@�����@�2{p��I��(��Pkϥ�D)�������=X�$��{����d�D[-a�/�^ތV�Ö>	�XS��˩;�DE&ƀ/��R���gB��yp�X��ƃ��"i��r��Uj���c @�4raϊ��[�\d8&:���"�C��L��j��3�R�}�G:,��S��?�j��y���}���'�e��!��_�m=��f����ڱD
%�>w�+c�c47ȏt,N�IbH(l�ٲ����r��-w,`}i�2_�P5��k�]���0�襬���$��� N{�hqx�+Ag���~�X����`1�� ������|���sph�pR��U�"?�꒞����jB�_�.�ʚ�+I=T�D;sl|D�3��Y�v	�/t�i�ݒ��n�U#D�o�S�Q�/���E��a��U���/]P5�"��BY��M"Q!]�N�������m�c%�W�D#��A��ʬ�ї���4z.3��X́�0��b�<�� ��Q5֕���5>�N�a37�r� SkIOU���Hą|�@�+�ᾎ�^����^TR[?Q����H�Y��@���&�G���:��:.� >���'Ԉ�U������+�n{�:��aEٻr��`qMI����VQx
�O��!��|�J��:'<�)s�5�Ԩ%Ԙ�{��X��pr2���@۹cV��+'J֍�Ot��HpEt��t���7�2FG@�S8q�Q�y�z-m\��ssP�wQ�:�K"4 ee=�E���V~�c���}<���C=�"E5�n�:_��lrZ{zx��
,�A3������Lz)E�݌J6������wz��S{��v��'�&S����x��Ŵ�����W4����P�A���:3ǲѯB��0%�Af�2��u�7@�L��,S���g�DD�>� M���I���rt#V��з؇�~;O�,b7j����
'p��Ж���X^QD�4�`
�]�2�z&���ޡ�d�q�n�z(/.^<ĥƝ��<���[������t��3�t���h��u�&=:9�'�->Ĝ���^Jt�`%q�o��B�7'��E;8���%�l5]�,dF�MwD�x����h�=~�'�C�$�U~�
߆?/!�0��_�DŻl�B��v�r�0���`�kQ%�;B���kś�dA�9�6����DV6揶k2��{]}�'+����?ʏK[gN�b'�?�hx�ZK���׊�~k���}�XC���ͅg�l���
Y��iq�t�w���y�)Тp�J'<k�eq��#�\LG�ӴP��#��k�r��fY��v\~�	�$�d���E�y�ʀ'��t�<��!�y<�J"�N�Π�+�4�~��0��\,���[7� ;��� ڠd���q���"7����Q�5ذﳟǑ���5��|g|���B�o��ۇ��y������H�*ϕ\��_���l	>>��葅��y�_�?z�dK�fE(����@d�U٤1�4���������x�����������Eo��g��ӻ��BB�z�y�Xa*���,�R���aq�6�u�����]AO�~��;��ChO��3Dp��)W�i�#�+5z�W�b<��=��*!�=9��!'TFܰs�jHm#�/�;n��>�A*�g����_� gQ�~�VOM�С�m��]�]4��#(a�K}98�k#�Z��9=�ߠ"�c0�#u�:8�И(9=�D��*Cu�W�Ŧ��1��l��/겈������H�A#�z���=���?,����B'�*���H�l���KK��N݇���a4��kb�הl3��Ʒ����~E�d{I�&"<��J3Ɉ�n���A�a�Dw�?']�J*yǇ\eE�ф���x�V��������NjF���Ʀ��  �v�Eu�k�!����Yҙ������ ��!J��z�pb��=k�;�u����nd�����ǈ�i}��x��_���em�D`J�+�E���2d��_ ��E�g��VF.j�̣OCF��)�0��w7� �\<``�4�I��W�b�\v'��vQ�PY��4���@1|�j݈>W�`�KE��
�:,K��
�e�Wo\ۊ�c��dy)$Y^�Hra�w���-�u6�T�>���^6�R�����^�i�"h󶣤'��z�ݲ!%��$dɝ���&��X�nk�u��U�����K�w���=�����h,�p�n�BnFdu�Y(����F�k9-l~�a�Ұ�[әq�v�(�t���M{��d�6���/�Y{rVN�拝ќx����~���1��M�In)����&ʝfc�N��J�l�vSd <�����9d��\^�Xͬ�\?AL��Ϝ�Hd�B8���Z�T�ԩ駣E0;�9�o�=\7"qOG�_����o��G<�A�`���Z�ʊ\��$vV��@R����ց��-n1�:U��"�v�I�[V���}!v�Z�[�n�Q���41���nX*ÍK۞�ނ/n2r�%X�)=����2d�Oi*z��ךf/f���-�o=
���6XbYY�ō��;<,B��R��-B_���Ziw�s;T9�����6�j�s�^�+���Y��W8��,}
R����Ůp�� �\��jy�u��fl���H(�}����LÞG�NzT�N	�	��c)�B��?�k�wR�F絯�d.�#ޜ2Y|M`Gƹ� �ٌrҫ%~@��^L7�y�<0Jֲ��%ջv�0��ֶ���eV=�Z� �	�5� Ѿg��M�i�0G��w7�<�,K���H�|����/-S�ު�*�3���+��j�ʞ����д��Yҭ;��2H;��Q���J��F8���S��~���<&G+�g:�H�gӘ["kI�qK�]�(^,IS��e|O-�֯�i]<�F��3i��6U�)J#��zti��G���g���u��r-���q� �����O¶�'jS�t�;���A���k�O���̤�z|��nYfh�cv�#�n���rDډ���6��v�������a����:wj���N�����P��ݞ�ZA���g��/�8�<����m�̾`� $ҷ�*��ќ%tl�51�+2֮V����E{t��ð=2��a+�1���<��b��{t���J<1/9/�7�["���#H������|�J4�ZL��h��ݹ�+���ܱZM��#��}����	��T�E�x��)e6
S��
D7Ylڗz�c�ӻ�'��xʮ�&�:��P[�]���y�TE�q ݭ��ׁ������\�S�J$�}�Qȅ<s��	 &l3Y��4�e(98��̩���*0&��ǔ�����@bb@Q$�F޷���s����f�Hw�T�c��g"�I���%t����z=w���C٦��q�y�}����4�����N�B>T>�E
U�~�ZR�_,�P\�m����G ��(V�i�q�96�3��>_�[.�v�yV>��yk��.�B�^l�%��[��y��#�X�Um�M,z2o��d;2*������p��1�������t?Ư~qҞ��,H���C3�o�c���}{�@�}�s!��_�&��ܚ���5.�s$E�� ���H"�����3�X*k�<�����E��w:v9��o+Gc4,48E���-�aGFr�q��#���Y�2Җ�J��O�3h���?j�'�`>�U�Yr��~F��۪ջMu�p屢��f�Nh��/c�tt���S=yB3Jrh��f��w~�y���p�p�I����p���*��yB�����kB���^=0��(#��
<K�V*i1��]{�R�
�J@��XhO|�[��h
������7M�i�+W���`f9$^��9�2�7I=j����n)�����;t��cG�K�Ro��e��+����i�4@ �ZE۫/�i�2��d_R�{��~i�v��ڢ8?�H�2���)�<�K��X.�g	ȷ�w��)-YO�-�
��y2ߡz=4���b�h.�/Z���ldO�ӜZ�a<B�"6�u�@�{lv)�g���+�%Xl�J��N���2[��%���Җt,_I2������K�|��ܳ(�����h�ye�dx,{��ޗ���.)��s�.�������z��0�Ã;f��zwl��Ҷ�~�4
-?���&�f)��-L�I�Baߪy��uh�v�]7��^�1�Kd�vM7����Q�)_�� 8�)��'���~���V���Ab1��/!��c5��2E]��@xp�x ���%8�py�0��%MN�(,��̍�TCǩ��}<$��1;cꇠ`Ng���^r�<�QI�"�舨t;FD&�������,1��c�>��	���{R��#W�P ,�R�P�K�����ИJʘ��%���$&c�|�Æ�V@#]��@Q�ȅ��c����x��elC#៣ �f�&��́ϡ��������c'�T��:�oJ�h:�8�<|���P#:ɽ�a	��w��Cݻ}�RM�1#��ީ��>2<�`Z��v���u?߸�`�&Ա-�L��p�64.�;�ƉL�i�O8{��J�縹���4ݓ��^�Y��1T���I�C�=��V2d���y����Α���{f_Y~���Aj�)��[�%�<L�Q�GOs�W���ٙ�gX���M��UxӁ���e9XeL������%������g.b�S�%� ^� I�n�y+�?PT�#���tiگh���4�DtI�$|^=��M/�%E��.jL�������I�bmQ"� Qgm4��^a�x ��E�J}�)]�a�4�&��SR=1��X4ھ��N�.�T�i�H~��л�X�/�ע�RD�g��st(M롃�`��)��4������� �s��F� ��M�L!��T�
{��e/��~���-����L��J�AB�ٶ�d�5�e�Q��Wb��З#�E��s˥%��5��	E��p�� ��4��_d��P��U�)����Ԯ��~C���MÎu�"�.�d��C�PT�����
�Q���pK��B]��`���C�'��E���-Q�0;��ðM�Н��.l�����|,�%��x"��)e��6�s>OD���l��:.�ol:�zWy3M����٦l�¦L6B8Ḩ|�M{�| 2�.�1?�*�+����2!��^I���QǼ��4,�lZ�~g0lk;7'rnQ��u;1b��`��︢��lR�^%�go�>��j�1��AO�׻�M�MybAXS��F&9�7�q?j�{��S>�+عk��Z�Ќc������N�E�~���OǏ�A��y|�ڸ�jR�~ƜK6 �<d#_� &-�Od��^���V��� @�����m��"���Z7<�s��I�7 �/������W��,C�A�8�M��Es�?;O�LWpL���8714W�m}$��fD)�$�SM5,VJ�}^��������vp�{���*p���:���>#}4;X�5F�t��9��y)�5)2Ķ�W��csߡ�[@�/��*+����+wl��:xcd�L3�av#�u��`�l��̤Y�&
����U]����Ӡ��t�|�f�k5��ܖ-p9�qP��d��/�X��y��qՠ��59�����JB0U}��ض�{�_�����F|`�2,6����4��xbyO~���N�ߍ��(8,�80m���Ѓ<�+����H�j]�>�\��^-���P�6�Y��<(���	�sr���΍9��#���L�U����[�����^�>�Pބ�b��[e��N]�*A�8m,L�	��Z.�S�dx��%u�%����WCcI����?+�r���<��y 4ij#� ���9IҎM��^4�������I�:����(�e䟘����Σ���F��R�6�|f�b�J�Se!���O���5�l���Eg�O������2? ��%y8rM�L$�8�P5�Z�g��yzd�E%ϻ�Q��rlS����W
]y	s�K\��ŵ�$!z���!,5HB���v��7g�E���C�{��� �?^�{?�zo͍z��d�B!��*͛��3QI��
L�1W��m�R/��^�˶����\��'g4W��QȾG�`#4w4��4iV\2��AnR�xS�i��Z��̧f�d�p��9ꐲ�}�,�f�3#4��E�3�1�;r��D�5�쯻Y��i��Ǟ�g՜J:
o��![�8^��>��Sʒ��T��?�#�������P�:ɗ�����M6$�9B]w�d6�����-슡;!g폪�!�=-�d/#1��Ȼ�o�A�ǚ�YS�����V襲�$��7��[�Gh	��O�.��Q_;��G�g��»솨���xu;�K�`��BV�]_���GL��:��?.�ո1 ���tU� �E	s޸3�/���
��֞��h�!u@��1Y�K�yi���E��K1`���t`9=Ú�[��:j������= ��(����E^&����Y�
G�|����X�x
�Ҏ���O�81~�1Z�l(���[]D� ���ځ�B�y%��I�Iȿ�>o��f��.qBP|8 ��=w3v����o|%��m
��m�]wڔ���4��w7v�H���e��g��_���{��`�}�D�ي+.� ��xUg���m7����Tu��:v�������m۪{O2�V�Rp��\y��*z��^�R���uz	r5�n��^:��ڑB+@G�X�m-o�g�C%��	��"kdV���acG�^�:�j�����+n�fG"T��Ngr��s�P����Z�Lt���E� �i�/8�m�Xl�<��5.(���HG��U���UݣG<��[ޞᵦ����Y�gIj����	��yS����J"�n(*pj�5��s?������pH�j�I��DH8��8�Wu�\&b�zah��U���\�a���{Y���'�y{裎lRq��kb��- 	1~�F�J�h��#T4�����b�wP�
2]�dr�}�r��mG��H�ٗ��d/猭���-[:ۡԃ���ث/������b���FQ�j����tp&�����EF��D:��R�%�l憜����"E�Ȅ�1h�+uV���4!B@1�DTi�1yVVf�E(�G:�����;�<?��B�3�K���b{R�j��nh��%?w�
e�����(_�U�BH�"�Z�b��@hw���mv9a���Ս����{l��G���ԞBd���e�k�Y��@�L�̓��s�:���]X_�QbŤ�{z��f_�a�~��~J��w%m�r�C^xF�8�n\���9��F���-x��O��pJЪ�R�ٍ��!��m]mIe$���(C��?����W5YOBV&����0�ȴ��ACGF��<Y�F�Gin`�#Fw{{���>ׇ7]�W����o9��Y���U�r|�6n�+�c�
 ����gU'�.+u�f��P(���o�{uEr� `u�+�3X��?�+�rxj�y�K��0H�e ��e���$c��eO�#�J.���L���:1��P7�g:@YH&�@�D�12̖N�&�'�S����z���t==Ǎp��B_�̓�_����@�E�Y}�.I��q�vCZ>*��o����
}�̵�0���͠T��fe#�����'ed��N�<	����7~ߊ�RP�������/O&�� �3�i'R;�G�G�Q�=���,t�����} �s�6�c�n���=+
0�9K��$�\0�w�[�E�Nw7���餈rDI����2����vM���|�:��X����
-�'e3�z�7XM����Q��W��߿����N4� D�H���4��ؼU�]���f�
I�-F����_�gf��Qh!g]v @Р~�C�@���5X�4M�6������"'�{ŝm�q��{b]UqbL�x|)+��>���������sCnP����"�^���"�ˏ��=��}�ӜO��M�@�� �⇰S�m|Rb`f	�`L���熂 �������Е��&�5�M�"G����r��l��wb�иB�T�19�9�s�����{��>�ΉB��G/��O�v\GA���٠ {�FZ���)�)җB_0(-7Ȯ�`5s�e�Y��;�LMz|Ъd��M5����sʖ�'=����X�/% �d3:�a�$��:�k���,$Ƶ���pUZ�Fyil������ނ<c�{���_�} � �T�s��I� ��e4УJ|<�Q�F�M���M(��C���/���O��
z�
��鶙�ef�k�z�AU���	N���y+KY��P��52��n���Z�I���;&sP�����jL��l��*���[��z#W���u(�JY��M��巜�������;�����+:w��/3���U��D�����ށ3�fG4���]���+'ˋ�^O%g|�i�SK\�9eu~�\�?dU�d2K��iZ��ˑ���9�f�$7�����H��wN����r�'��.R �6��'T��R ��ɿhgL����C�����߉��;v�0>�
v��Em��ög���/� ;��
-����>y[��Aէ�a-�����$��,���<�E@�:Q���)��2Z��kꜨ%N9-0����^�P���"%Y-���;�<�Vb�����]Ʒ��܂��}���X���YWѪ������Xvn-��ǣ�m��ӌ���v�L"Ql�eyD큥UQ��Wg�I.?���
P��X�"�>���SF�5"�Ah^H��!B�Y�₅5O�����3 ���\�Z9輅����,�)�G|�r+p4���'����%|WhY�`��Y���9��"��IX�rr�����V��Ҿ��ǝ�"�,�QL����ð�U p��nk"{��P�KNF�>H�b�s�������X�J����ɑ�D
����;4��ٮy_��/��X�<8P$� �����_��K�w�����eK�5���C`������W0��,y�X(Y�i_�>5�N�|�ʩ<�G�&�+U��gPԲĝ�]+�u��1CqƸ�l�9�R[_G.��3()�R@��p��K��RE/,��VB�#TnX0��@t|��9 4��� 7��(~ND��e̋IR3�dx����6b>K����,��L�X��*ץX��]+�+6CN'�z�/Pr�5E�ha1�4�����m�f�Լ����(�!�P1O�u٠���ި9���g8�I2_y�$1�ɀ���\����~å�:Ge������*�0;[�o7���V>��Z;��U�",B�n5�K�Ǫ��vn�DvԃIo48Bz�Mӱ쌭<}c��k���
7���T���ԋm��Vʧ�9͐�A�;��IP ��tM��P��p��]A�FU�`+k������ �3TAf�=`+o˗�/��ͷ��H��|�Q�w�t���J㕬	��n+$Ն��Z�w�j�;��o�u����	��f��|�ũd䦻s����l�F��VF~�#�k�����������%jT�,��ӄj���ˀ~}cm�`♹MrB�Ӥѩ��>�+^%���y#��D�Mj�+n��a�Q���Q�(�ϕm�g�#��~�[r&�<R���=A�f[�`����v��=�u�x��2�����2aۨ�x�@mc�+�s�A\-����2t&�p�"G��gR�	d���k:"a�7��2��Ն�8�������$G|��g2��/�K�*t�eMC�bK�P���(� p	�S7(��͝?<Kܫ'��U?�����9|� ��"�m���ے�!��4hʽ	�U]�$!ڎ��B1�X�X��J�EiU�X�_�X2d2���>AH�DV��k��Gl��h6އ*�����N�h�:��ʐ����s>�YH��9�ą�Y�������;�+��0�bRi���^���iǳ!�/Y)	8�_Ja����.ί��#��x��$7N����QQ�2��~��>�������.$���M#�q�Y�����G��7�BAR���\� \����r�V5�$���u�:�}��� ��Lʯ)��Q5pڇY�݇{Ô�)�yR�a�V�u>�T��ݬ8|�[�
�2�ӑkoؼO�#9m#и剝qW�+��r
%�^���Fb:�6���+�A)!�ktY0Z���!����׾F���:�"]9/ݟ����d����0�g�:0��-!���*�%g�]������o�nx6�D��r�r�ײX{��Y��h���?)'e�ײ:~u�la'ݠ�Q�Dg{��W�#6���)�![([��4ee#���m?�S�uq�W>�\�=��������!���{�vI���M��.Ԯ��=5��4������k _v��Ɛ��Bi����h�]ɂ*�¿I�K��s\���zg5#�%�W�*��O���� 1��fC����3��%�V����L��6$�x��/��`y����d�6�DQ� 𝑖O��-�܀"��_���p��i�cJ�Fa�AHL�>�E�T�揿���Y�ɀ����	̓�ꀂ�c_����;i,ox6c#vPa�2�N�75�nhmp�^�4��?ߴ�Z	�������XtV�uA���KS��ϭ��E@-3l���yK4�W���z�0v��f�\�w��B��g��	�����q��U��[�593�7J8�=��ˢ�I=
��-7�w��P��wN��g��W-��"�z`t8'�4`���IQJy<����^A'tȝ��
��H��j�f�x�rY��b�9{A�5�a鼈�:>$Y���8c�x����^/�+���kQ���TXk��ʲU.�N���
�Ǥ�t'�N+�ASw[�K1���j�a1'��	՟]���(�/��{	���'8j�%%�<m�>�s�?�f����۔<���A�=i.8܅�$N����٢�V���|�8&/m�~���.q��{,�7lS��Bn�4i"W�̙{����Aˆz�|ꋤG�q��s�j ��ðe]𻷐ѢU�N�Sl�)f�wĔQ�׫���+ź�DG���,��xU�=)������ҕ�]���y�_���2y`	����< �(�T�*��uvm������i�����ή,[T���A����(3b�K&(�G{��f� ~џʪ�,u��B�2%3��7�ZP��\���ĵ&�y�!�M����\@��_>^?mҵ���S`I��۩�;��ÅTI�ݱ����3H`V�B��3ne����g��#��Zǃ���;bm1��u^��
������)��F�#z�#��C�"�nx�oh�,���KL� 6�GG�Q�t�Y��5M��H9T��s���4�}+V��1��m`<�@�n/K������H
�@)g�y0х�M�No4I<�g�R�徭_��?���)�U��k����K��?AҝÀ0F��o�%O�Wۉ��m�#�����m^�����7�����BI4���1KP����I�(��>���f9AJJ5�'��=�@N�i(I��'��1u��1��w	�bܗ�S�+ϽV+�*���mmJ���j@��(T���(C2q��9�~q�c���]a`��{��*�˽d�%���Ѣ�+P�������,$�0p^Uo��ٲ�@	�v+&��1��M�E�3@6�6x��R���#-&�`~1C�6ڊG&����w���:�]/�&\_�M�p}!��Q,��EH���MVEEO߸�˯�#>������%�(y�r��|�cj�x�O��[�g�`R��FD�h]���p?D#��7���=��oO�S�i[P>Us%K(QP�i����FS���#N�M�bz/��W��K��.�SS�;jV٤$�C��p���
�����@G��������%fM=&-`rxu�Q�Z��&Fv�:�UKR�Ȑ̲���(%�C��Sg���w>�ȏ��;�����CQ=�>�R��N��J2|�L��v7�X�����`�=	8V�y�;p7+c�0�V���m�G@��;���h0�m?ΜJV�~�6^�T�)]no�֪��/[�%���'��l��a�[��)?-���'��>��K�S�j��������dnyo���m�)��m���8�tDEĸ��k'(&C�-�"��g�ƢUl�
�̧��9��#����kp��8�Ih��!*��]����2�`6n4�ȳ�<"�J'�'G��s'���n��~����hF��t ��v��%��t����j[���6���+�w��Q� ��}�y~�h?u�8�`��//(�X ���ͼ������%m�=�-�M3������ro��<���,�5��zLvj�w�a]��S��%��ख�����8���P�6�5
P��y����Q⟓g���(��g�x�\}*R|�}@�?|�ޥ�z��0����n
$�` H�zuw���Hh[��ђ��z��(���;�g�F�,o.W�&�rK���kJ{sM_�䐫���(�|$ǟ(W��0��衁mc>�x��~��;���v��Di%^���p˾���,��e���q�"g�{�lb	% �۪���#T��S/��sX���A�pՅ��=��`�����c���VDG�<�	M�֣���w�K�2�Z(%��FȄ��v�
�R/b:�CAQ����TU��`�x�a%����&��ł�ں�0J���!���5�<�����+��0�>�Z���Ro�#؂)�TY�n!\0@�A�x��l�#�j}�e���U�eP���"jl�`����)5oW�ś��KS�4>Y%R1S��,��=���QB#�/>���; ٜ(]�C
��D'��6{3&�(UQ��`B��o
����s�͔�I�:k,��a9�Ѓ��K��h͜X������p��xj�x�u���R��tc�sX��d��%�C�\e� �U.��A&�R�lyܮ��7MP�ʴх��Qi~�9�7��ٍ�o��C%��&1�	G����{�,����b�٧Ā�ܽ4Ii�[�$#e�;�"�K�H�_PJ�࿭�BZp�c�m{n��2m�N��n� �@� ����RTFT4��í�����ñ'V
���]�,��8+5�Ɲ������rg��sp�&"�([8M<���k�nV���SH*�
Q�鎢6.�f���DU7�� ��=�,N �?�T���"��O�,��7�y����D��o��H?��S�k	tc�}��rW��%Z�A9�`�F ԫ�&�!c����$A�����&8N�{�v�>�l��#�˰�� �j&Ͳ�0{B���&5�I?������3�ߪ��3�dS�8���N����,O3�A��>����,�&�����k�xf�*�I�sy���ݥ�F~�e�P���u��al�{��"5�������̴Tz��{4�v:�)Xj*mpF�e��m�ݜ��I,,�=�E�2̟8���C���j���n�}U�^�U �lt[m)"��ϔ�2�ty�4ȿ�s���:�Ӱ�e�/_`$_�0�p.%
#�/OR9!�.�;a$omjE~%��7�U��SF��Q�w�/fbR�ZC�r������[��!��l��K��o�]�
�ǯ�2�6<��
�X�;��9�5��#J���B��>���T�:m�qJ�(3Z�`VO� �f/�/U@�=D۩��P�O*D�Y���[���х�Ǎ�k-��TĠDz��1��2&n�۟�V�� ����B p��r���?��|.�w��{4���P�AN1�|�e�` H��,?t�W;��'��A�M���]l=`4�Z��żs�������x�X�