��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su˸Y��'��d�Ay~�`�i���o3 1&����1\T�����	��!mF��
��\�ݘ�#X4|'�~a	N�1�""rϗ��?���ݝ��^��lt����d�k>O@�0�#/���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>	��l_����b�-V+�t$������b���Uّ������)�J�ܮp���'.9�|�ַ����������N����E^��q��;�`�[�`��A`�?���%J^\�N�%�p��>ER	��.<��M�@��͘]�-j����r��O��'E&�_A��lߴ,@��+"b�
O��Ѳ�m���ҙtM,yĥ�f	�𘶼0�'�����n.��Rs�l|��Kcy���a,�r�^D��K�1��o!A��Ҕ�BZ�� �ؗ�ٕ�tצ�|��)8�<��%6 љ8���@�/�w�u�(bĆW���ک��,
�-02f���rs`av�=�Y�w`8=��g�	<@L�9_���J�(��Q��nU�v���@'����G~S�D����\U�1�����������)�><��-Ul�a�V%�Q�j�����vE��>�qC�M�v�`ym�G\���T����# 1l��'��"�E� � w��P[m��#`��'�7��:v1^��!�����{�� ���~�V�)����W� ��C�W�����n�c�x؊C����U�'T�h���w6{�����#2 ޻��F�|M�z����<� �}Ed@{���w��qI9t}��-	�S�N��M|*V63�_lxUUTx.��	��M>�Y�>������{�ZytPy<W0���"��}�0y.�i:+̦L�`8%i�[E1�lT���^��ZԿ4��`�4��j��J��I�N�.#
��΍�+iR�+��~C����Q�ݻ}ü�({T֐2�|������sPJ�+��%����+�U=r����4i��6������5N��� Ef!�v�'���E��en
(a����)uP�ESB��dD�M5�فx�@����G���Ǌ�^Jzz�k;�ȁΕP�\���+H���ZEkFZ�Ks����������d�>Δp���4��9	�t`eq���c�d�%D\E,B%��4�#ʦ +>��_ɛ^������̔��CU�Xݲ����P��r���q�(b��CVN�ך�v�~X���Ue�f舜�h��=�A�9V��^�����t|}Z��I��P���2d�u5�'��Z嵼r��r��h�7#���4%8�� �o���� Ow�&|$����2�a\G1�+�q�
�}�'rڜPL�뉫�������B��o=FR��c�Jk�ݍ��4����OgC|�������4�q��[+����bn3��T2��}����2�B��q9pM7t���� ��x���M���W�F���b�CD��ӅҜ�?�A�ٳ�d��\Y$łmI�����n�-�3��cb:���ݏ���2�f0����z!t2�?q	w���[����5�/ոm鸲>I�����/��Ͼ��í��(j�%^��@{�.h��NC�W˼���y�HB�4�
�	x�,��o��<��`ƿ!�|w�H�o�72���ţ����T=Β~�Ш��u6��4����׍&:���5L�g�[����������}��@�3�2c?:�;�]>�B���,\�B�Ch5^�%[���^���j�/խ�.ɻ�8x`��%�����3iy5N�5����f�^�b�4��G0l�2�,�x����k^w�]V�xk(7q�=�Ɗض�(�Xn�Ԩ�C&�l8Ir�bW�V������/:/��=��c���o��@��Wc=|�(�
�I"��B�$�a>Z;���ӭ��6�' �S�ި�=�����
�F�&����ԯ��0�)O(ga�'o��;"̉K�z�.����MPG�'�����g��rP�Q�(%�Q���������?����=���Ik�L/n��S�R寕��ߙ�<�K��e�o��&c\|\�[Vd��|��\�����z��Imu�]�ta���s����uJs#�����I��x�ʫ���,�ٯ@��ܦ,��X�4�����A�E8f����f+��q�c��K���aN:X��^d�SwI؈����{��qf�O����*���)���_R��]�y�
���G'"���sԨa���>{��=q��$	�g��	����~>��ݭ(:�+�ފz���A�A1�������h�Ɔ΄��)�(m/<�C��J{n�b�Os#�)LY�g�F�8h�εZLQ�+�����D4�>�R�N�P�[�1��"��@��k�z�7�o2���)�lM#�#g&3���4z�O����s�$�(ʝ���ei^:Pq��]��9���[�ۯ*:k�᜗���;�u�f�':$���n9Ộ_L���I���y��&�Nee��+���N�?�;=,�r��O��!�gsX��{���i ��8Z ��H�A��> Y�L��_�Z�X�	�4=Z-���Q�g9�{�)=o���<��Z�$���mm.K@d+#�<�J&Ȫ�����)��"X��q\��s��\IO��S�PC?IϢ�eH�*7�F����R��fs��3d�l�)��82;�O��j��z)�j�Z����ԫ3������?R,�ؚ����=W�7I�įx�[v�ę�o��O~�l�².���Gع^��4� DW§�Dw�9>�o�)
޴
}�� ��'�4���sR�<R=�W���B?�`&.r�� ���+��*��o�D�Z���qO'�����h���=�#��Ӧ��,,��}�Z��1᳀�����~�rd�``���eF��k���?�F�(�"H2��9�^�|o�pw.��VEo�Q�6� � ��k۔��V"���\��u�W#v8jh����Zhc�|c_��<&�t�z��P�K˭��:n|�����k��O��5�h䁪�?`l�d�b��9l�0���\�^'���~:X��u�w��bY�+�%��iEM�� ��6�T�ٙ�^W �g׏n;nx�}�GYcX�*��E����"�n��G��ۜ�_��^_��IB���k�Xc�M\��G�>O����dْ���~,���88ҦB���L*�8�,�C���tX���L�(���"C�:[Z[Rƹ2��� b��`qM,�Ǖɴ���g����EMY�imEr%>�'7&�yp�{���b���K��ED�˷��iiޜ��FPx���=���X��_A�@�i��W�,*�e$ �1�/�JdA�����OgTI>Ѩ����Kw�*�������9��	�]h�އ@lh?ֆ��?d������<��x��`dG X$a�v$�>��v���J�&� O��a$��y�	y$#+p9f*u�qا]�[�� W��C��^�|}�P���"v=3����^��b1*d����jY�eK�ʣ�20%��
�?N�s�}��cSm#d'�z��Nm	>(��� ����.o�	��
�EE�����G�j����j?��ԕk��t���^�BU1Hӗ��%d�T����L����
�LಝK��L���Z�\Jg�I��[*��F��1����+�q�M��Er_�qf�ʒM~�/�Z��NG`QMF�\��V_�#�Cuk b�+�:�%�lL3���?��}c|�X'��y��]���ʢAת�"�{57��[�퐎hQ�M��L�'D�ٜ<}�pe����,�m HH�٫+!÷ڽ�r��ie���`�����ͧ����bЋ4�=�R�%�wڋ���>x4���E�ѾNt�}y�K>�2����"�3v�1��OOv	1����>��yT�Z���򇾸E�Oȿ�42���G�?5z4�5xt��m�7�*��P2��������V�%ɘT�wTJn�.�~���T\^����-C8c��ea��Q]N�śj\;������3lK�-�o鱔@߄�	a����S/Y���豿���y�6�,2v� �3n� ���Y$�[0�FKd�m�*��4���0{�-��+�U���dj{�@��e�f�#��NV����4ۀz�D���o\�DcUm�&R�T�	��0SXu�"��y+�R|O�Z�+���"���V�(����)�a����K�Qu�D��������C� �?mw������$��f��=\p���S�c��<vc-�q������ف����&�ڷ<����r.H'B^��VJ53Z�U�`�2�/)�����~���^$2�E������G؁a�s�@">��`Y��ʩ��]t��7�L��Dz����y!������$(�+�����ꪯ���/�����
��{��Jt�;`;9n ��>)���b���<IV71"���?׏lf�u�'��Ջ$¦b���ʌ8�/Aǅ^����1��J�eEA�i�'��cc�5���z��тK��l�jTVf11���pC�Ya}N�����R���3\]�P�P�v��ѫ����@����t��g�lt}��lP�o����vQN�ָ����