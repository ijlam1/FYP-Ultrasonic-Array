��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su˸Y��'��d�Ay~�`�i���o3 1&����1\T�����	��!mF��
��\�ݘ�#X4|'�~a	N�1�""rϗ��?���ݝ��^��lt����d�k>O@�0�#/���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>� 0�ʪ��O�;`��Z0`U�Z��	aI���gt�3۩��g�Ze���T0�8o{��
y�����%(�3qt��M@��w��sé� ��}P�jl+o���
���;���^ =?M��@���^D����5�9N#���wľ��l����Сw�c��FK�JH��O�<���퉟�
�=@N�_\�p�_�vN	n���S��MU��T���O�S��y��x��ڋ���x����-ӣ��9}��-�SZ �b� �P��6�:Q8N�)�-~H��ڄ��ؤ _��f����~�����E&�C��W@RQ�ݫI+G���ي�mgX�C'Y��CN&�@�ʛs�W��0֞�D!ݟ�a�ߨC��+��D�p��nq&~l5�.�<��7��2��y��w��43�hn>�̵��E%>�x�p�uǑR��.��?�2tU<��6�N#Y��r�w���r�Sm�惀�C����W� ����mL�����^>��eA��R�~^���øu�3���֗q�:{?'S��ѾQ��=Y2�
���&�]^�,C<1�jXw�ֈ�ۢ�	��q$�H*�7���#��3��]��x${!J�%���IPܺF�.]������E���U�Y}�������|G��`]4��+m�F�D���\�X�*F�Q	�W���%wN���u&҈VflK{�f��o��&�G��9��A�iBQ�x�NG�J��^ן,�@1h�5A���'�-1Kz��d?�U���ǲx�J����e7wZцA�9ج��u����	3sVR�[�ӓ�\��hr�N�\"�}i���D��qx�3'A�	�$'ٷ'��|�1֨v���|��!���wB����M�A�:|��e�H����[��뱦���3��g����R�#J��a�'�j��PJ���E��L��W���ƮC �&���ϩ�e͚H���-���eC6�KW��`浒���v{��"���:s��;){/ģ<�W� ,��t�C8����`�P�c�\�O*����E����lx��~�<�3@��M�c&rʖ�˿�ya�J�Ɗ��C&ײƃH���8�ĂE�BZV{�|p9=*R�t���.s!ʸ��x!dR�C�� ����S6t�W/�F'O ������.C%����*��߰�d��j'��ans'�U�e���r�<a�k�����"�W�m�(S�8�|߸����Ӓ��s�l�d��#<�+R�1_i��_Jc�"��j �r�|tF`��U��ȶ&�h,i:<~٧�42��]��~2UAY�j*�Tom�J��n�FҒMn��]�z6��:���,���q�0���̈��b.rН⤄#��9�� Hd��X�s���
m!k��e�����j���I����$Zt��ITL{��(�.z�Xǚ]�}��RFF2%�|�.m�զ�Ij\GZ�=.35Ф߬Ӑ���E����6�0���h��7�*��� �]{��z��5�C�%{��-�ly�5�R�Q��p/�x���t����E�G:�~�П$���A��
V��X2,�
�v�w���ۋ2�[37���eJ�̮h� ,c��k�#a5�ԵD?�������<�D��!��JF^��mr�o��W��	߸�+wh��= O�ǆ�y������3�Ԧ]�7"A�@+���QvM���̬���p�2;��ꤙ�S�Z5@�Ϩq��UU��K����Q��טɟ�8��Q6c����Z<�m鑇8@��[_;����+)3*;ҹχqX�'ɐZ��)�Wʾ���aw�S�8d�'�m�QtYTx��֞�h>�빽Å�����tS��2�yi�ڇ�#)Q�r�}��!��� b"6���?�}t�.�}H�D�dB�[2͑.���6�6�~[�YvXD�J�!�ņp�Q���?:$Ke�E$���J��o�1��������ეX���'�#�d��\��	M�F~�-�Bq3uj5�f�Y��ZBG���pIwgf���w����v�a�&�~;��x�R�E�iU>�}��(�sl����Ẕes�v���`G|�)K3瞩�S��}'`����q���SU'����n鳆q2�2��Z��8�܊�/~L�L�~$/$w��}%��X���&wα�'�C�~}���U��b�H���&��vD�c+��I��Uf��*�nۨr�JZ�G�~�7Zdy��L~�mދz�϶���W.���*�Õ��zi�A��l���x^Oʈ�¾?)|�8U����	h�5��)Cߎ�x~�J�:WTR�D]X���@���I��m���\]�����Y0�qk�|B+�	��v�a
~�v`4�n�L���ޗ�l�*�d�U�Ǟ�n.Pؾ�*Ơ]��u�w�=蓞����ߞ����N6�ȫ���)5�������xT2;�Wb;��F!:��J/_���G,"hcݐh��!CK��ɏ*��� �\z &W�)���7�Ri10-U$(KB��;�O�(cbRvd������1Y��VT�S&��U�)���73�u���C�o�um1�.�Ƽ�Ÿ)��.3�zo�b���ݵ�?�p�AQ���3w�����<���U�%w�'X��ަ��,&t$�����h�BY��ؼ�?����s��NV�[�5�μ���,I���L�=�C>I����C���b3��崶f��¬�7���A7�k��}p����߮>$�Aڢ�	�Ⱦ?[U�qFr8_"jk�qz+��"/��W��`������×��Ώ�+�Q�}�� 	v��dE"�熪���Ú�ДV���Dr�*��?���4� f�Y�f����5^�8���Ӟ�M�۳)�mO��=-.�u̱�&�/��T9�+V��*d49SG�<0�&!GT�D31z�H��P$�dlm9��OK��4��ƐCD[Ҹl����'�|&`ʀ���4�4���YK����ye��h����6�ib $7xl���31�����/
�5�2���՚$�1�Cϗy9g^�3j�q�0cW.)+�03�T4�Q�G��4��ޝ���kK"N�1�������_��LQr�pn�%PQ{i�z��љ��ћ�06�8's�1)�4;L�!�>J�4��Vdi�[�{!42�E�#
�>B]PJ��Y4B ��H���_�qj�$�Ə!�Җ,Ѻo�iD&�y7V�w�pha�;�Ҷ*\ca�h]��)	�6Y<ԖX�"�B��r�A��],���kPw@�r� �<���K��a8�	E��q�e���<����J�8z}����v�Q��ׇGK���x���ض�hN�H����'�l�2A67�Z5p���$|Ȫ����A�}���C� ۯQ�˲��{t�*�����uux-�]藚��̶U��_��"Ʃ�