��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su˸Y��'��d�Ay~�`�i���o3 1&����1\T�����	��!mF��
��\�ݘ�#X4|'�~a	N�1�""rϗ��?���ݝ��^��lt����d�k>O@�0�#/���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc��3@���;��̵*T���që �|c\
��`P��o]L̛�鿕Z[<eLl˭�W?�;���Xo����^����Z�<�F�g\CT���/4�Ǎ�@�����(�Lx)�EF}��N�QÑ�*�����Zf�ϏJV�E������V�M>؆1"��0}��{�ƽ�`G�%[�,s���>�ӹ*����ںA��j�'j��''$���F�Sy�,�v��i^ٜ��/f���.�n���WG_�kQ
-,�.UI��ۉ;��Y��ULCͷ�,lY{
��B���<�����N�CĖ�Y���3r�����M�Y����M��<S���K��p�.t�<5���EY�Ӈ֋A�3@E&%z��)�܌&ѹ��	���,�6�WR���D���4��QW��O�Rb�9���5��3z��Ia��󯏎Gj*��m���1�#=�S9`|�|�8���F��Cٸf�;+�AP��{�@�PT�����t(�7�wg]�����(	�;��S�f�W�m�t�x;f���൬X���3�p��r��9_��Pή3���}��R��u2"~Za��nB��8�f9���f��;���El�Ī)�a��J��m�o͛+̒��P�5k�N\/�^�V6�Ġ���>hO�)�cɫ�A"�N�Yb��k��G�t����_ѫ+� �T���c���ymx-ϼ�j�~u��y���e:-�1G��hK��v���@���"sf�i��Ċf�XB{�����]~�=��ϥL 4��-�AtCFSg�z��j�%<��|1�,G� ���E��bPp�j{��<�"��R����P�
|��m�^�/�~ஞр�o��%�6�jb���N5c��T��򗒛p'�C��$���"�eV��<��kڑ�	Gպ(m�� �;>�f�1�B%/����������L�wF#�V����q0J=����8:�@rP1�N$�1����]����K���0�m����+�~W��!�>��,�ZU�>�@�N�Â�T���� ̱�Vѷ8�j7���P+o9i����-��``�2agk]��U�}�Smd_�7����-@�Z�	N�] .ي�h�s|֎�����3�?�kxx9�J�Tﱡ��i��nB�j0�>{R���9��x}��&/H:��+�/���d�;	H�������%kzr�����W��h���i���ˡ��NK'
F�T�}w�0��b�[��a7�M�oUh��-�&lP�z<uA+�]��d�\�&��Yt���Վ�P5�YQ��$>��S[c	�6��k�``3]��]�h��&�Fӿ0@��Q���"eGL��.0h�Z�OL|8�I��(��i?D��s���
MpZ׬R?�Ϲ�R��{M(N���Pe̽n����CQ(涷�r�E�9q�o���������9�>a	4��}uLUM!����g�|Ã�;5<����@Q��,��9`�iN���V�����+�'N��=���q��H� �:�O���*�wqy�����I���&�����ʓX��������q��d�`P�!mO�r6���,^���T���"Ԥ��\��8�Xb���o^([�h@O�O9)�k��m1v�f�K��!Ɖ����ܶ���M0�H� �������l���U|�������zF�^���5�-H��G9ڻq��`��D�h�O蝿����� 2�B'c������w"�"��J��ߚ�<��:��M��%��+P�]fi;2eF,1h�&���F� y�K�F�?գ"�1;q5��U'�|�iF�(�^/ȾvY-��B�O��n
�3H�Z�@�M�#��_�Ԣ@N3	)�V=ȶ|�FhO%�Z8��H�(oE�Y
d^�[@"��R���OSϟ��30�MYIH)�R}��3���4����9���D^��j�sj8<�_�;�ã~O���3�0�
ӄ3ƃ�<5|Ѐ_X�� ��4z[ܼw��ߢJ�mq�V�J�J0R5���.�_1Id�.�X����~%�|k���,���;η=���4���KJMC��c��%�y�=�H!Q��RC�K8m%M���U'�W���Z��}���I�p�����܃�b��Z�{b�fޔ&�Xu��_({���Z;_��6m;Lɳ��8��̵|�%L��j@58��x��ٿ�Vic{�q�OC!��n�3F���u©O�xr�_y�8c�P���{��Vv���T^݌!��}��Q耓�|��"����u����C�?WU�ٺ�j�Ӿ�&�3�n��0>���S�6����[\֥����4X��v��i5��1PC��N_�6��ɨ"��ތ��-�ôz�/�:�e��n������sӆ)%!܇m)k��4:��v|`��)� |�wK���l�ܭ�ǖp�ǭ -�SٽW��g���9�2H�-�X�bg��>�F��|}M	�d��O�y&�@EiTW�9�����G蕲s���+jS-�1�$`�V�';M֟��3��������3�LG�
�ȗy^dn�lrqp�9�LJ�k��_����fƺ���+x�kZ.|����1D�ؠ��v_%$�-�ն^��}9*P�c��Mo>A&�U�\����&<�)������[��g5x-���5O��[�\e�u�F��on���`�Ne���B���Q'4\`�
=�9���)h	������R.��r�ee,�;ǩ�^4��;��Z�b�V�u�sy���:�Ѵ�N���S� X�I���IE�nT[ØuXǝ⇊�((�@����"�/���S�D* �<�<.~��L��Q����)Ujٔ��Y�ۚ|���wT~<��&Ӣ4�1�*�j7�[�Q��a�@*�����|!�s�3�e5�I��"r0���ŉ�Td�W!��(�
��j_�f� �p�F*+-Q�^�U8�.x