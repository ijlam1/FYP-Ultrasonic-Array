��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su˸Y��'��d�Ay~�`�i���o3 1&����1\T�����	��!mF��
��\�ݘ�#X4|'�~a	N�1�""rϗ��?���ݝ��^��lt����d�k>O@�0�#/���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htd�X�C�[���0DR���a���k&|��p^�GU$)˻r����f�/V,��[���e�k�ϓ��)����y���/ul����tތ�<��4Yj�[�T=��� <e����^Gͻ��N�/�]r�|�T���ѯr��=��g�]!��,IRo�_�7�O���'&��m��@�c.:�D�����GW���B�n�E^�_�}��d�#&j3��"�J�����K�ߟ}��II��
g�P^Pp�����'Z2���?p��<w�P��#]��"[�
'�q?�E+���t��=MJw��$�5ٍV�5�0�� a0z&��<m�sHU��ZMNq�=�1Cpd�(�u��;:M���T�8��i�Bctq�WTQz7P����eۘ�����I�u��.t�r/�d	�%���IlΌ�H_"Jn\DUtR~��ۍ��84�/DS�(v�q���5�/���5�CA��4�6^�V<xC�����%'x�e�e�=5�������a~�������cr���fO]\'� �_��/ZV&j�nd���S��Wf�=���|V���=�K�	�8��1�� d�쪈�	}�?N�Be`����%�gI� (��x\�p褉�5n�4mu��$&�l�]+�S:�*o��/��>������d���u��V�����i�	Gн���GnMKy�cD�NxǏ0���V�s 3��'n�St��t�lQ�������Щ×1r��n|;�L�K�ܪ�y���n�ҧ���u��_�`|^��C�[�Kϴ�w�����y"�C�"MX�1�9V~�p�#� \���P��X�(*�+=�5�u�U�Xu��0d����*r�p~�`���*B���C)�5��C��H\�#.&.��1l�1��O�:j�r,��);�ޑ�`�ϧ]D�,E��ϻIP+{�=(��)A%��tl�d�N�3�r�}zP2 �Q9�3�K�����l+ˎ�Q@F��H�|���I�,տհ2FKW�f�9��컒�%&�����4򲸋�����c!@Y܆f �S,	��e"��T�r<�dïvD.	!h(e�Kmڨ����~���|d��3�e�Qb�9��zf��;������h��=].F%[xDg�H��AN!��#b3���dh���ՌcU)x��z�B�ʊ�A8#�*70��V�<qP��ʛ������"!��I�����I��02��_���<P��]~��;).�ƒM��T�m����'�<�)��P�z��a�[�?iKR;��?+ (Dc
t۽�K�����:���'���y���6+��c�v?�B���
jS�D)렇o��ŷ��m�	n���ˋ��^T����!�Ť{u9�{V�)ӣ���i+���ɬA�n>�
�\�4����Ҁ4a�q���}~��oR*��q*��$B
du=f=�u���(GH!㉼���=���m^�d&����S�~ ,JXc<��e���� 	\�������	������#֫y����\�vy!�C��#�t�V(d�ei�����8�H��7T�J��rd`'ϳ���l��i��U&|XUj����O���Ǽ�{�fE��%�KaG��5��L�fp��m����C7g�z5�B7�R	�H�_=U[X�Լ'�qX!4����u[=8(���w��R�B�"#3]K�y������Pz��o"I+���jT�{A G�[C���6Cz�ӟ�.j�M;h���s�!�r�*���( �r��r����냜JW�Asb|��^*�9��H�C.v'����Z
q�:S,1�k=�a��34y���u�� ��q��[���Ѥ^Ym�PB��DZ0�x��6Z���l~���3jcb�DJ\	�b�=s���Fi�Ff�F�d@�U�#;B8� �� r�ԁh_Bn���s�����Gx)���ޠK��X ������8`����t�a�j�"+r�U�y��<��������2�Vs4jŒ�9�I4'�	So���NhΦ��p������hq�W�(�}�M�M�-J��z��y��ͱ�^RT恦�S���Y�/�#Ht 4�M泑�V<R4��0aRB�\m����\R�-^�0��T�����m(4>R���l��(�3����yno�m9κ����F���(/��B#el��1>��CZ��IX���,�,��
"�:��g�$��yx�����9�B�iYi��K��96�pMbh0n<�g�>�U�r��E�����Tc#������~�ӱ�aw}�B�VL��TB�l�"F0W�HO(�_���sD#����Y�\!�\[��϶*�,�y���
=��D�,,�<��/�d.Y���Vģ6�2����j�j"3���*��)tb��;76׽� ����Ǟ+&���$�Ѵ���������*�|�_pP�S%?Q���#0��={n�����*��B3D!k/�U�f�j�(��7�ch��8�Wɛ3�8`ߌ�u�ʈ��y(���[���Z����J�T�1;Zk�z%-(s�H�b�Z����'��f7 ����g���"�B#�'&ķ�[��%�Ԏoģ���<��y����m�!,P��G^mm*T£}���M?��?�S����� �B�����J���"a�s�%���ǂxZ�&����2L�P͟�O՘�&�9_�%y>����f�(쁁{~}�1�Z��>Ʀ��D
��΢�ŮE9���)�g*Q%AF*M��8N���2~O6���`�]H�����¸M�ԑ�x'�2_�.���D}�E�`Ԗ�mO5Τ�)̯I������<�-��`Hc��t���k�r ����8��K��h���g����U��D�L��<V��ab!ENc_�7pj����`%Xc�%�vk����Ih��X���^0p��OU��Ȩ���Z�p)M��Pzqk�����즌���#�;�_N7�r�I��{L��m�zS0��\Q���d�Q�p}`�t?B�����n=_�=ǘ�S9?�AލF>�	3!�:P���yu	i�\Uw��<���5\�R���!�U�miu-!�V"��7�&U����I�ě5ì�<�޲����GJ�VBV�q
!vNs��5�PՐ��1��Ͻ;�������I�5�_X��r�g�Vٮ���~�v%M����H6AIL*�փ" U�5��~ͣ�[ ���-sd9f��q�@�#�뼱�������1&I�!I������b���͍P��-�\$o��;1�Τ���/�(�JP�݃ONyag��sAee��^�Io=I7���b��/� ð�cB(��̣��A�/��guZ��
�