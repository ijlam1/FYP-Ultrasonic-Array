��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su˸Y��'��d�Ay~�`�i���o3 1&����1\T�����	��!mF��
��\�ݘ�#X4|'�~a	N�1�""rϗ��?���ݝ��^��lt����d�k>O@�0�#/���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>b��z�PP k��R������֌��pT�B��Rh,�f&`?}���<F�Lr�WB� �Yg�Rm^M���������^Ā��|�!�!TOX-��Č�Σ��z�L�R�;��I��G(�����-v�*u@/%0z�1�.=X��P�i�~KdN�)C\B8��_Ë��uъ��tM���#8�b��3�`��>�C�h���`i��$Q�x2S<Z���"�o�n#C�k���1_�G伨�������N�px�L:���CQ?��OU0
��$zҀg��pm`� ��]�G��}2[���4���z�ڥly�7�@k�2:�#"X��C���6�#u��E���=ȱڛ�re6~ԍ�`6>_��a���4gW�,_�����t�b�Fm���/�HPb��3T�붛7RIFtS�V�r����$��-�j�.�8,�=z�g�� ��xÏ�N���^O�(�ADgλ�W�[��4��o�⮢n.���\�	^�zD���Lh:�X��,�ܨ�A,d�+$�l��{������v��?!�6�(u��`%�SN6s�S~?F�on�kq���y��FBס�M��`t�h��+y^z+_k.�p�X�;Zb|5��m,]��cL�t�)
��1���3�I���"��!K�B���Ҙ��컯s�w�N�Y�T<�C۽����Xk��le�k��4���9:I�Xs9�J7�+�а 
�X��|t�m�9�-�_ݟ��R��N�`z�&�>��^�媄|���n����JaMr��T��}f���%^DT��]�G,�G����5�A[%�Xg!��[��Oa�,�vL��)����*I<z�>������N?�d�?�"����;2���Ι�;�?����b%%��F୯�	���ÿ�ʗ�l|u�Zf�����)��:���w4� �'(� �々��d�g�8�TX�_�WlMn��<�3?������r���D���׽U�W��<u��h��`�^��@a�)�W�Y�A�&�@<����Ȃ���~��~�����AS�(��9�d�͓�Fm������Y�ˊ�"~�~<� 0�����s�>��OJ�|r��2TL���
�Oju�<+-]j"B�쬈Y�V����z�2˾�u�X	�4�E<H� 6�R�֎�j��iǁ��
�3W��i]�JTs�%��W�ZJ��K#��k-���ҙ}-���s?�Ǧ*�֛�؞�%r:m��GU�?����]�@q�	�Tˍ|�݆�U���"��zV��.z�v�Q�&�M�&���_O�z�rT�j������+���c�;�6'I���7c^㠡l>�IWB<^D>�F�0��'�x��3�[<Ύ�-�?j�?�v�&��L�NV�R��!��������x��\��ɪ��n���|�>�t�Jq&�L.�	�;��\��5����yM�3�5'h�cjx�o��p��t���׵R�`�f�x/[E>9yE���5����x�x����]�v)��]�Y7�댯���L�FT�0��7(J�@�~)�����L
	�������o����M�q�̕!&:ʇ�y.�j5~��gto0?�C��LK<6�F#Jk��U9j�����0E��8U�ق�r`�J�o|�$�}^j�9��;��hf�-���0�24Y�O,�C=6|E��k^b������Q�W���!��� 7�
0���~�=Z�s�������Z!�𔒬F��X��y�y!_"I�]w���v]�?F<�pk�>_�hQ���ۈ�_�-!t2�m8y�F����2	`1���D4�P``���S�>$2{$���G(Đ9�x����B����x�(��2d��O�b,�]�^ H��"��:Cy+�{ϩE��%��>J>{���2��c��(h���G/�eJ�C2@cqfalI��l��1�^z��7i��b@vg1��5bnH�9�I::y@�.������,mw��]��g
p��W&�}�6�%��ݚĔq��N��g0���s�&4�U:>*(����#f�͏mL=�Y6�`�HS�7��y#e�:qa���ň Ws�+[:i���הI�\������e܏�֐��
�a>��B*~��u_�`�\��i�}0��¥B���}]C��f�*���ߘ(� l{���Y<qʊ��
!J�	Hd���\����O����#Nx�	�U[��~%��l�Mk�តG�3�Z���� zx|���z��pX�o!@����c��q�8�*D�]z[���Hoav�f��чFU?�UG�a�5e�8Y" �x���A��ԭ�J#U��&҅��9T����([�a�i��'���G%$г�hÂ�-@�x~f�S_^�c�}jq�;N�i�at��}�$���+1��|��-�����.����ܵ�:-~;sï���0���������d�Ѯ�Ue��a8���w�wJ�l�VU�8D����a$h����|�ߜ�#�`����h�K�����Q�����˖$�bJQ^����R���?9ԉ�+1���{�QNݘ����)���?��6����9s0�V�6��OG����r�1/�TK�;�=���|�ڨG��2R�x8X$�{鮕T�����
�T�$�3���ξ��C��ʖ�Юk�1���L����ٸU���H$"�A��Ex�ZŬѸ������}4�ĕ=^��X�����/hh��?T��N�X �'N=��OB�@6��B��E?]m����Rh�P���`}K���6y����Μ�u+P�=�������e���km`+��)��v���bQ�E_��M�K�:�Ty��Љ~��}�~����;��[Yo_�f�q�k�ŖV6'����1k�:"%�ED��7���|��YNOB@���Ώ�J���b$v�y@�s�C>���+|*��r�6�a��m M �KXb��@9\�{5�1;�pS	���QdW�y�Kծ�H)��è"�6y�5I����]�{�����aa$D����v�>��k�aËD�c�Gxt�k4by~у�L� �}�YsP��J�y�A�`o�rre%��s�Q��u� �E�;��a�zJ�jc�>uU���Ǎ�@/2���|j�Ɛ�}1��|� ��_��]l��nw�
��d�.��&�0�d�!<5VM3㽕
 upa�o�i��#0�/�dԳ����^�EdAU�1T(���
���Of��Y�`3m&��X�ؾ���<�nG����)�����q����D�~*��>G�
���H]��(������兮\Q��Յv�p���J;���)le%`I�By	�:�E�˰
j�����UT��i�3ÖJ�^�'b�������*	�[�|8�
Nf�Kʟ�\ofY���%	�g���bCnrF/�-Y��p��H����Kpq�D�XRV^g<5�<$B�b�?4��q9���"�6��!!)d�E�TcTt�v�-����OB�JYd����S~�
X�E���@V�n~�*���E��͠�ٓ�X�Ɉ�Ï�~/)�C�>�E[[A�3~���7"���e �d��5�v�Ku� �5 #;����ko�pWOx��ox�.���څ�Y ��N)���m�~��A/2кd��U8��d��'"��m�^?�.D��1��(��L��vrC�l�_&5I([�"��o�䴯^lt��Bj�%�TA�f�c���gp@��C

�C'���l�prR�h@k�vh�'e:���Ś�LOw�bU����2��l	��j����&��0�	�h /.�G�k@��/'��"�z+�lh��_-�� +b�Y�=���Vj�M1��.���i��0�'@i��/U9"�cfsc�>��K�9k����/0�o�#��,���Y�P�	H�fj6s��0߁Q3�<�m'��P�`jÁ�`�;/|yp�!�vH���o'�X�B6?7�k��W���?	��u<\�k��M���x���	�� L�ML��ԗ�����z|�Ń\�-�mTOs%k����>FDV�6ݏb9�yp�ٯ�q_�D70�/�t�ŸP��L���C��A�z���sa=ׂ�[�'M��S3 �N�D�ٵa�]��iI��dE��@��ԃ�v�:MK`v	k<#��_:t�	�4��'�I�*dkX7�;�#�G�ˏ#�����30k�a�k~NX|��[0<D����W 4�N�d1����-1G�"�49B�y�a�b�MV7D��3�#�1�����ͯ�|yD��a��A�j褎͟������l��0dg�����`9]J�+Z�����\/�\�
�mEMM'h�yI�����Z����7��߁���2�Ή��M����G�n��p^J(76��>�7�U�M�z2bo�aRk"��'�h`�1�K�� �+J�\��WP{#=3qаI�y�$���o����x�
e��Y�0@@�`/9u���p�8(؂�0��y�'hS����l�'�T.�]aSzq�9�'Es�IЭ����r�/�w_��P(�W32�.z�����s6���p���9��ڊja(�\��W�qL���T~�D�q�̏gY���f�\�6���U �$0�ʘuC_=�n�V�։��P'���Y^�< M{���Կ8�[�s�\��}I;If0�1��~Ǥ���P�STd���s��Ǌ7! ���(ޘ s�ㅓ����K��N<���^́�B����&S���5�JG��®�R�I1���.�bP�3YHΉ�1��F@ZC���_�Lk���r�zp���g��h�~��q5��v��,kDA��C=:{C�MJ�_�T]3�I[%�8����� ��Ē�Ɂ����K��^�cisi��0�x&�)�I_��iwM���'�f$��l����̕��߃�� �-ςz�.�G����h7)k�fF�~��f�m����
�4�`JF�oԿ�m����\pK��PȘ�xO�K����kRՇ�Aʷ.�?%��� ,FD>󠛟���BiA~�̭�����0`�-�摣 ��|�e��4U����:�¹�Q��;���zE�|�`l$���.��Q�UbV���^� Q&6�!b�)v�`�$��C�t',^����!3I�ғѐ}?q�?�:�FJ�݉���Ǿ�촽�Ǟ,�����qY~r���n,��������#�P���+��f�C3�,Ӌ�l6�[E�6�b�#8�X���΢&K�@��c_yh^E=ȱ��:x�)�@����f+���h�y�(�! |o�g��뻜���ĖV��h����)급����'�D4�h�h/zU�f�Mn:����n$�O�#[�m���؝-�@c�S-t0�E"�F�%�֓�,�f����ub:j 9L��2�#&Mc�x�`�-,w�qs�`^����߆���"����jr^+qj|�D�F����AZ|�������Ĳ`�r�B�=d��-�$_XQ�:f�F�����y��zK �`���-�9ѣ2�ʽ�8����fDl:ZK�-�6�����+ћ��	��gR��|p3�;�y�o2H�OKZd޸��Gc�r����(#�/�~M�cp��ʄ&��x�!�O�t&�c��Sm��~�z�S�3�G���'���<��b�e}*t.�IeFՃUv��SQ�øFlT}�����_-�������e�N���~sb���$�{jn�܊ z���/9 �q8��'|����W��l�(�/7G��f�C�#vtµ+C����HW^H��X����/��lTVȉ�r�����J$z�C5f;���"=y"3�.�\3h�;k����}O��,�$����~��;Т��?��K�yђvc�U���:K���z����㡖Ŵ�%�C�gzW�ю�����ĕM#[e�dYz����@��Ƚp��y��7Q�!s� �c�}:��MI* ����t|����%v�a-�j�h��x"�����k����A�W���6�GD�^8�[8�ho�<q�r0�����e� �T�FZd��z�Ӭ�n.=���J����$�4e"��n�5���)�H����$m<��������F��g��ǲ���h�6���x��vy�%����bL��د^�Χ��,k �zʠp�N�������~9�_C��������jo�UrE�g!;�h
����k��@��,�u^af_��8#$C��� W��2?;P(>9��Z�U��w�"����T`���ưJ��vK�M��2>�Q�}���b  ���P1N7�γ�$H���dG ��M#W�7�Ң^��[|�14��U��G��e�a
�[R/L��Xe�y9�X�����,�aѩ��S��OW�h�,�