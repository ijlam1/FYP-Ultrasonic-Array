��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su˸Y��'��d�Ay~�`�i���o3 1&����1\T�����	��!mF��
��\�ݘ�#X4|'�~a	N�1�""rϗ��?���ݝ��^��lt����d�k>O@�0�#/���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�7ټm�lQ�חY���Y�IW��M|�O?9��)����U�F�\P���qm-�ň^E� ��C;c���6��ר��QV]P�x�u�Q���-��Xҏ�R���b+]���e�	��j��7l �����ާϸ]�y,�����2�<���<����q��f&w�ů|�23v�8.��l��kw�KM�2yNȇ��u�&@;:�Z���ըq �x���*���l	v��k.��������8���CNb�f2�������z���-@�V���(�x���/�e�v�w(��iI �cS�g�c�Ѝ��%����x�{X}��y�aZ�//e�1ю��UJ!��D]�.D���Y���}>�1|9���c��?��L��4�R��~��%C/��~�y����h����Zy.-��D����j���E��0WhY澑�pSp��%Yy����>�q�[�HK����,�[�r�)m�2�G/�@g���-����}��7T��O�� (��O^j��*G�ϟ^!�����_����#�.�ͪ)�ǿM���Xݦ�p)EQZA�r���'��!�ß��� 80&G
�%4�k
n$M�o#��ڣ�y���{��XO8��u_�T1`��fч�Y�y㑪�K$&\�_�\я����� T�_Oy�×z
�q_u�Z� *�ZP�i��ON���� ��螧̧�C�0���Ƃ6&~�b����k����M����
�Y����on�E�
��Z�mtP���"��!��l��y_�����z$e�K���\m�=A�`m�\���1�m��͋
�L��8*����A����nt �.�n���9(�kb���8��a�޺���5�G�^3�"��d�5o��4��"M��ww$���D�,s�����v�^��u����NRzt�[_n��rL�Z��g��T�V��M�`�nZ�t��w>V��B*f�'雼��)�YVה0�AV�XN Ͱ<Y�k:����;����ݝ���1L��ْ�A�1�E�wmx�����E$񮐧�so�͉�ڇ����5�>��*� �*�����bQ���_|�<�q�Zy-d|R�~O4����܃��wsy�g�;������F����%��qJ+��-o}��ݝ��iQk�]�F��[���g.��Ѧ�dMy�"	�1�$���6�ζ�ʩ�6c:�w$x���V�"h~G؁$x �%�ï�)��[뭲�̹瓱K��\�c/E_�>[F"�J>ԧ7`fO�ǖla��6���g��sۿ��s��;��v�����m�{m�clh�e$Ǜ9��	΅;�2顿�������UT�iJ�df��ޮd7n�݇/�Iy�d�m�lu;�NҌ�w�7��y�UxA��U�/��T�ĝ� ���N6�,a�Z�(�z������F�g� }�A���2S>סr�U�| ��0Vfኲ�,���a��!śO}��?�v�s���?n��ݧ�N�_-�b;2��a<K�g���Mʀ*�R^ilQn����٣��"�M��E���D[LN�Y�]-\Q��l�-=��@
��[��QQkŘB�I�����-���Y�a��Nu��Wc�$����v��x�@7s6��X��V��,������Z_��w������ʜ��x�=o)Ƈ�	��a-y��}�2�������KC\��:�?���ΜT'P��~��T>p�Ц�hO�j�܁�"%���|���4-�ݹ� U�.��1��UO��F�����1�a>�B��|����	�j�E��������9=�X�HY��_��;��E��5ǐ�	�K���p}~�5	U��w���Y���AcI0�#������:@j_9�liwF��EgM������d��Z��#��2KF���Kjv��>֜�2�~,4��Z;�,�X~�v_�Z�����ae:�<x�6G�I[�b�>%�7]�Y��\�2,D��4��W!3@:[�[�&�h��Î��cN�9� �ɮ�P��Z�<��u������O��.����&g�䙶q�}��S�]��pq/ۮ���r�!�،P9�(�BWFA� �dK��!L��I��W �%J���wF�B�|G"ǧ��q�͑�����[A��7L��I�Y�d�a��	[z�%ʽ2�ޣ	��G6��K�&��g}tCV<�� óo|��t��1�b���b��9����9��YTp1ޗh�>5=����.Rڇ��F�Ӽ���8��Z5V�c���n�~�߃��W�ݲT���6�C;�&G��g�Ҕ���aM�r��D��zo�ٝ\��2\�����?�P�h|&摑�1��-��v�DF��c�����9�\hL9�B�<�a����p�n`�/�F���]�ɾ��J2�6e��ڤ��N5�� i'[�c��>���.��1�`ay���k�C��qq�&������B�Q���B]�D)ɜ�2�'�Z���i�jS�����z=�n�F>�U��>��t���_![�N�e��bF�Ƃ	�)=ZB��l�Ϗ�&�T����kW�?]c8&�<�ڤ&����%]1����7�➐��Gh"��/q7�2�0��L~Jfc8���{���G�
	/c��L �L1p������Pj�����eg��z�*sL����՜�/������N��5�햟����#���N{qt���⃐1��X��JrMT1 f�L#%{r�u��y�kO���Y�lBu�k$�x7�Z��ΑG���Ɯ@j���_��L%7�)Q+D�c�<¥���>�a��8dmA��j@�r��;��[�q*е��t҃կ���
��]�_��`�h��h�	�'��Z)�b�M�JNm�wg����S�.�zD���ڈ�<�&��؉^6�V̄�{w�fsz!v�