��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su˸Y��'��d�Ay~�`�i���o3 1&����1\T�����	��!mF��
��\�ݘ�#X4|'�~a	N�1�""rϗ��?���ݝ��^��lt����d�k>O@�0�#/���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>���q�;�;�g�?�_�q�-�m��5ʞ�œT����
��cFZ��R:�'��o�xE[�I�N���B0ˀ�2|:{4�C[�p6~��n�?�Ϳ����^:٘�!,�i�dF��<<���0������� �Z�=+C�r�.3]rܕ�u��׼��)t�C�n76�ˡ��Ƅ����;�lG_��es|V|M�m��=�^�d��F]A5=�M(�x�O�y���jIAdrg����ӋiS�]&$�c����	��5��6F}���1�IK�������JMY�vmh��@iz�S�����IjY���B]��6e�?��X�b�Z�/���q���v��ѻ��]���TJ\�v�*ǅL^�h*n>�D�[��Unǒ�nQG���+���	kD��p��!10V��m��:u<�_I�e��c�,��h6ʚ"��;�_]���)���Z�H�2nz����+�G�!��2��Q���\��wa��
ҔQ5]���X`k�A��#Ƈ|���P7R=lN����m'8١$�߳"��'��.Y��!d��LB�,"����K	`����TN���:Kp��C�Բ>#Ŏ��8��[��YA1��@����\GOz��G�V2mŏ�W�g������O���L_t��W���[�tQ,]�z%����_^������p� u��+�Mk����Vr����)9�� ̇nLJW5}s���Ԩ�0eb:b�X�zC����cM�û��+i&�������s�}�)7T?���Y���A�$GϬL\�QuI��,/���PX�'N��d�-V���r��
�WL��.!
Jo*�R�e�T!�r�K��6��/�.�$F�ԁ���)��r��P@�$��$@�'��u���kɯ�#�蹭G�U��u��-�?O[�o{wPb�N��[^턃XT�7�T���)Y��������M�QX�K��x�s/��u�͎�����o��w���PO#�%'�#����Vz��߹����^��E/zV���_K5�`N�k���=���V��F�Pi�NJ+���|ӑ6�2�o�ο]��(���oq���KX����wn ·��Γ��7�K�s�����+BK���h�PFĂ���U���c���D#D�+JW�P̆$��-߳��p!�Gn�N���я
G�c�|�xTq�8��Z�b����> �[�bv>�g�<tEL?xȽ*���N4Zm���jv6�W�x͊T���� �K��FM/ASkUꥒ��dy� U9�UT�FJ���)p\�Vh����Fy�9H��LR�k@Ŝ�!j���b�z�K*+	nnG�%��1��"�\{�q����Te;@Ϋ�9o�UZ0{ ���S�H���HT˧��6����D�AA����y� ����Q�4M>$czN�y-�<u��I�����从V?n��ĵ_F�ӑ�L���+B��Gn�IX+��~�����?m�(B��$|�DC
in�h+_��� S�bDu&��p��:����{�R!�UT+�Iυ����~V��j�Dg�RC?J�� }3�`�jh�����'|⢱����׼�r��W40Vq+=��U���O"9_,��E�F����)�n�I�=��+5HT�Y��E}J�2��} ҞS��e�ʙ���`/L��C������m�'7Q�=����V�1�kKA$���˕��g��L�I���@�R8�'���Sx�D�2R�Z�/Ȇ�ˢף�7���S�fҦb��zV Œ��V���S���!{�o:�{�M�u*��s���B~���2�؇$��V�3����	%!LD�����f�S�-m��ǧ��<#��b�n���6��9X�I�$\-�g���?��17d}�|�G�(� *0���+�%��,�Yt�r��E��!f9"9�9M�%*�1 ]{g)Z'�X`at�CK�1꨿}���h7�\R���@q��={��F�"c�q��<�*&7���jb�c[l��E���kM<?g���8|"����L�:G�N��m������vl�)�l;��{����.�R���%���8�M�_�n������${ D�{�6��TR�cpm;L��`���%�Ͱ��
��F- G݅��O/-n\��>���� ���Ƞ��������/g��w��H��w?�.�^�2/O�!l�����{�0]7����������HC�>=߷��mI�g"l+��җ>W.�>�8��sOj�[m��V�̣`��`{����,I>s�#�^Y	�ذ_r�@y�&1s����,hP5yA�A�Ӯ$?@�O�BG�%H~/T��;�ZF�l�>l2D���$�Z�stÝ�m�1��Z�4RD4���GL�[�,v�����2�8uߋ��Xp,A[0�����PO5�$��E�2���6s4���o�'O��.a8��D&/_b���M*D=J1k�6�͂,�k,\�Ia#��4B ��Z�aj;G�XK�w���#��h��o�a4�U �J(�߶��@")b��^�0m:M�J��5le]5������k��3������^
�ցw�/���j%��*�EƌV�٫gү���R*�m�|����∭}�ʘ6��]��hxՑL��0f현M�K�rX�B�������0
n�`�`��\���uo�L�r������;��Y�3�IP�PBBa�	`qi_ ��huBu�C0�.�-D׼�v�I���/��p��e=����S��wj��6���G��m��Ò[��	�W��޽�\5��c�P6�{�p�ua�����ME�x�'-�|����5�����HO��ϵ<�HLЌNy��o7;t��ud�9o!�}k�%3��4�x�F9Ho��D�0s�P��; ���N�9�dӯ�9>�٤�o��&�a�9)��O	��L�6��Hl�̐֟)NX�Q�` ,̠�����֌�����.H�C�'�<shy+�tV���1�4��� p�x�^$�S���!��N�9�J�����-G�q������hJ��O�e����E��=�R��:vLU�h��ɪq����g�0�_Y�`ϒ���]9"��'m�;'R�|$)�૵��� x�0OT��➯��7zؒ��^GN`!���0�s���Eʨ�S����azM��_�����g.�n�V���P~Ȱy:���ѷ�L�s��ļ5�쿶"_3b�I���_fߐ4���G����F�d������{F6I
Q�:�i?v�-�(h*��8W�?����wI������0�7.�oU�Gf��;B>���ٝ���,@��[�Tc�2]��ĥ0F6(�&�ë��g��/j�F����<~a��{�Ŗ��*=����XJy^��Bߝ�;w��!�,�EѼ�Q�#!���v����j/���*!�c�+��Y�(���������<;kf��߸�`��V\�w�6.��h�*$���T�y��55য়�����1�&�\����@�K==�;o~+	�EG9�)�#޻�SK\��sv��ΰ^(�c8��X��qm���%���+m#��
5�47`�}�D�O�[y<�����E�����Z/��mU��J��[B�4�Y�,.*�*Y�i$�G>�Z�;���H<�͐���z��8�I]c��n2��!���u@tW��[�JU~rA���d�1�Ԭ�w��29le�SS���u�,m�YV[!Ô����҃��#&?H��3��C�5f�i»��Vv�ۧ�D�/��7�dfZg�=���=k)���<�L, �'�2�N5/�x�Λy_j�K�>��]�ygAW�e9堏sȼ�rS�R��z���!�(\�Ä��	���U�؇�j
-�������e⚢�(Q�.���n����v{noh�
/6��5M<�l?,mn���Ljd{�����E�y��Bpϼ����7�"<�;���x����A����!��?k��I�e-�o��.A"e%�9�Dl�1n�t�\��Xd*ÇI&��C�,��/	���ch������)�
�ｊ��v�M���	�#�X�QL�M�Z̤uNH�?n�Ȑ���o,�E*G\GY-��Mf�=����}��M-���%tt�Y��Ml�Ye�_!&���K:���݈�~�I���P�7m�ۆdf�Nr�lE&�ˬ��$��\�����R��y���Ri|�������8�����O�օ��m0��*'�?�8>NP2�̶Î7&F^jk��������~�\kǼ<F[%��63ա��Ƣ��1~�j���sXݹ.[V�(x����Ǫ������X2�~c����4{#z]G�ٻ�$���xBL`�4�τ�Q�ro��*�&��Q�C%:UMF#8z✲�Ube��c�s��y0�o��e4�q���B�.]��3
��i����lJ�W6h
�śB�QtZ;NN�^Q�"+����k��߮����ʇ�M
��[/wSZ1�R>��ա�dx�^��3cs�\At\\M���u��s��Q��Bڱ9���2��H}���Cϭ�C�g��#l_W<����]�V;���xc�z�W<|�z�G���9|R����>�����'�x�� �hg��$�;�����6_��H�z��*��������������Qy���zǂ|X4*�}}0�O��^����4�"y������%M�i��S]W��&�^mp�\��r�ӆ���/�l_k��	)#�=މ l�G�B�C��G�Z�0�Q�E2��U��.a���~�0��f�W��w�#Pg�#�	�\{�@�)��r,Hc�%�%+���J��q�/�
�1�����Io���)�ka�/me�K�[����8.�7�t�9�a�5I���M�a��@m闯�MA�$W��f1�L�7jy�{�u��$I���P�O0��
�%'<��v��,':��.�q���(�~GA�Ms� �V�?�m'C6������c�1�lQ�;;��q6��-|�utFg��W��i�W���%�3�C	�Hv�x�xt�	����I���cO&Y6���_h������g�u�i�T�ŏ�B	Y$5*���}8Z�Q(em6HT��x�q���o�ʵq�j��^E_a�v�e��G�:(���t��L�9��Cl$B��B���B)�X7w (+��}ۢn�;����ޥ�z���Q����Rtl��b�I�����g�K�0�ek��6;җr@L"����m�-M�(��:^}��Oum#c2DSw�1�^:�:�AN�s[+�JV-�A.�V�l��VD���4�?�9/��F����Qή�ڒ�"���2aŴ�ew
]�Y����ƜN���Ns��ʒ�*Y<�έ��r���5���ym�A�ɸ��0�X��Դr�/�ĒX������]3�<T�j+t�i���'�Cx�
��a���L��0���I�|�Ӳ����Vyj��7Ӯ\��ڒ�N~V���;:�<֣��@�:��8Va����_]��'�@r��|�%�"+-�����=�+AUY�I@ Ϲ�����n��t@UL��ð���{sj�o徊h��.s*`��";�Zd$�Ъ�ff��ݽ�mY"��.����f��"8F�3.�v@�Ɠ>�5���s�l$�
Ǭ ��@�s��@��A{�3�}���̼�%df[�ދ�q�:.:�<���s�����s %fQ6
X�0۱�S�1��]���e�>
�U�c�"Eʪ��d�wT�(7M��H�5���u[RU)���qN�/GK�{�|��S���M�t��d�R�ݙ�ײ�><l�	.uz�w�rc�y������}R&��4�b�0B�d�O�AY�s���$���?w�!��JL��Y��OIxa��/��SĚz��-s\R�T�]���� �ٱX�*>Ա�*�u�����U6�J�;� �I���P&��H:���xsi37n�Yi�/F���/9s�$e<�1 �ub�Rg^Fy�R�� �"�#���/$}L� ��h�Mad�$�i��.Moo���y�a�,�~�R�a�wꑃ��{D���y˞��b����e���u|�Ki7,zƏ_Z=8�(Vw��	���s뺔U�93QzU�<!��v���l��H��Ly��q(�K��1g��!��i	jf�#�%��>#�m���+��'���3��]+*�ҹ0$X��0Ov��cm�ĚA��EYUs��`�<�Y7�&�҇���6��e��m)le �����P�Ө[�HzGG8���?�9�Vk��d;�8��SM5���E���X�ݶ(���ʯF��)��YX�2Q���0��,Gs��(�:"z�w��|~d�Gr҆�Q 7RW�yѱg���P�˔�Lk�ު��=J=�,.#�+��=�뺸ð��M#r#�P�2�/6��_��:"��k���hNA�DɄ�4��"hWd���G�� }�Ę�a�b�<F ���R�x	�+<�`�J�h�fk��I�TS�:Q��h��G�;�Y������l��#m������.���1Tطb/��G�ma���M���:�4i�7�v��CZ�Arj����/��1�O � Ķp"�F/p�*�r����җ&�>�P���� ��Y��W���,�c��eDcE����	mjn��9�̶�ȉ����ù�+2�Tk<P�J�ܨT�o�E��/�g1l�ef���kn���0�d���0�íWK
PK���h�ݜ�/�#�SQ�{N��O�Rx�a�Dc�4�N�����P`��� ����x�A���(�U!�_��7���l����gw��l.�f��+'���\�y�]��<���2%6��[j1^��E�E�-�ݮG�W�̄S��A�ڻ�^�}����G��qt����V������aZ�h�"d8r���I�"_��\w��5�9b�`Ƨ��>9�������1��5z��ߨ<Y�f��j�*�,G��	�T�\t��n�2�툮���1�J�s.��mz��b�.vs؏�G����h��/�f��\C�� �����Um�!
M��H��R'���Ab,��?X(�d��n�g���v�\��X_�V[���}���^�USc��>|A�Y �J�w�B��N"."��64����]"c�ǟ�#Cǎ7����I����Q�.�ϛ�*�b<�u~�f��E�̽�X`��v��z��U���ڶ�Q��F-�M��MO�x��2Ϗ�R�L"pr�"1U�(i�����;�4n��^ȯ>�"�ͳ��#� �>�^:����2��=��8'�ԕ�c-�+v񤄢��a{�Hg�����I�|3~|3X�~\Y��j�N��L{�8O��bh����c�NS��ׄ�Nn�ٟa���z�j���;or�y���]����U���i���b���>�X�	JΦ�Z)1~`��QZ�����%O��z(�ԣ��w�ԋ�s��#�ٖj�pc�X�*K)Z7K�f�G��_�c�xh�|]�üU*x=)]�l��P�����p��g)�'9#��cy��Fx``ؼ�q�/{ ��UC:�?����#����[�	lG�^K�RKfɒ��9�|�I�u��{Ҥ����n�������z���s�����?����,-��9�Z�r�џ������*N��p7 �7l�h�"�:����z?I�'����5Z�m gLz�߱��l4�Q%����F��b7X�6�n)S���R=���
u��<�d��^-s�~ʏM�j�ݒF��f˧�q��n��{���u��3�L�b��8��ȗgsl�o�������@�z�y}�Qd*<~�NK�!�[���0!��Ȋ~VLw	�Ȗۗ���M�`�oFd�EFKK識F�"R�f�d�{��y1`BPrfY�H �~����X�p��|#*pMw��|���ԷN�_#�旽D�.�AH���⧎\�aL�.������Nc.T���v2Pf3��EKԈ��p�ȵI��8��Dc�SN�d;���6KORO��0	RK��_8����K���{A���3�_�M� ������l���]ѕ����J�r+բ����1Q�w>�%~�;a���Ӈ�E@/��Tb��Li~�\f��H���D=�r��\���e���w䠆֌��.So��\�"U����'%�_K�^���R&���c�������!��a[�ef	�96�b�$�ĖV+�m�33�J�m$0H!ne:��&�f����Y|	�/��N��gW1��z�����4sق��Q�mj�Y�^�6?������A���	�g+��m��>��^��������-C\_��|<�I>�=�a�3hu
ωy � IkOLf?���D�m��n�X�ne�ͼK��zwH˲�<\?Z5�m�_�Kp�I[� e0��>�S;���m�F9��5mh*\_�b{-��3
�/�'�_�q�I�v$p��۲Dߠ�[
'�}(-<�e�g0�?3:�zn��l3�C����L�[tp�����.'��O�-G�DۃS뜪i�o�12��XZ&j�r\��w��k*�G����z톘�W�qJ��u�a1�?�5Ds��X��W	O>��ed�t���K7��R�� �N��HWq�%w7#,�)��Ǎ��2����轄qb��HՑY_���6���k�	BOlS:� _��[��q:��W�+G�"���F��v1����NN�>�L$h��wO߱�Zs�ǳ�o-H`؄	��p��z����������c@$�q51<���u�եxإ��yt���.�3V[�x���q���[����V<��x�,�2&d���V��3!e�r�q.�"��m����+�y����H���2�@"{� ���@gk��1�	�ƇT�_���Z�}��aL0n����Կ�wz��_�p������"��@^1�ya��Hl�v�0��~+Yu±�_\��H��ь|��`kk�o-8V�جC�c��n�C)��T�ԯ҈�2!�x]�u��OQ��^�8�i����G�csm���73Rg�$��b���*�c��!��P��$b��tw��Y����2e�W�Ɉ���A��XІ2Hŭy�`����b��>_��,���+�ٜ���ztQ���ѷ�-[�޷V;��o.��kF����%Tx?�t`�5X.ѐNH���r�a<0>ׇ*"s#�9��|`��P��{�ߌ�(M�|�^෭����b]W<o��lW/+��KR�M\]�`$tE)Ɋ~��APf6�&�G&9g̰�
P��yn=�Κq��L��e���gYL���R�;CC'b�-T6�f��yA�}��E�H<xɵ+�2�[4��g[��	�懲_=���X���~w�y�W%��ɳU	��C��c�@��^?���Q��äBqهE�F�kjG�Ci�[��8�S�'<�<ж:b	��m��v�ŗ�Yj��疓�@��羂#����	Kj�
���a�,lgj�������xX���k �o�jK�=�N��7��M�����˿��ɓ��ڸ2-t]fqI�J�ݨ)\�|� t~f���F����~���!������cK�C���ov���^Po[��[i�/ � �@��)l��.��=�68�5g�Dߗ���v쏋eP#��'�Gn�)�\Ep����ع���4��-�c S��ȝ�/�<I��MM�lC�3)�G�U�3\�i_P�9}����ǃp�U\0?��Z;�ӷ9��*�&��G�`݄N�F��S.�b��f�Nd�P��C?$j��^^����7M���j{��*,'�#jS�V=���Ϯz	[��S�+!K�T�br=�z�+��M��R��7oI�$���S�*\�;?8�@ݘtڠے4��&��j��� ű�� /�:�5�ڂ�A��nd>"�_���?j�������+k�����u���e�|����N��T�o]`�7quހ[O�9]Pi^��&N��a�n�b�o� 4K@P��/{��jo`u�W������!.b�
_��:_K/��>.�B����W�m�S��yZ��_��3Y�b<������ro����'w���=�7�\�o]���Ey���lFe��r`���w0�f��J�g}��݂��ur�b0`��Z���#/���dBl�[�d�s̜۷�jNz	o�&���y: ��o7~�9wT���9=i� �"�7��g4P��ԾA=�`y��!yPA0�kPM��8���+z!�;��O��U��$��-R����[�{��%��zs�����j�s�Ó�,f@���CIS�'�d/�K�]�~���pce��h�Ԅgi?c��#ҡ���g�^����dt���\q<�w�-����\�
�"�����dK�W���8~�bU�7�0��)V���l	������/�tN�7X۰�;�[��'7���`J �d���pedA|�k�5Y/�ھ����;b;��"*�c#����&&���Bx����IA�5+:�6��M�9hz��NɗtA��H̞��*owj(�|�=m|�*������,��{�@���>��t�<,����S��I7y� �B�L�klwqKA��hw�2���ϥoud�tH'/$oD#�Z U��L�bΈx�~��֮��#���ҋq��#Ɔ��F?u1���66T�a�G�YB�N����z�S#F>gݏ 7H?�:49`.��1���NԸ�̨
�nN�����J6�X��&c�	�M����(�_��b��>&X�~g5\������M���.a��}a���~@Y{nK�~�F/J���Rֈ���G�څ�X��K�8BZѱ>^��]�e7��c�b0*|��������,��a$5��sQ�ڊ�ˤ�^��#+4ɺ��xK{z<��Pz1i*����fN��U<$2C�Yϩxh�D��@�l����Ca��G����t�{.!C3�b&�T�l��c:yg5e�qb&�,#�<@p��bb��3�*�^� �OG	-hT͊�r�� 8h�n��.��<{�'���h�^~�3!)��Ye+�Z����Ju�]��:$I񐸙��i\� j���f�/C[�/�)��׃��������"U���u���܌����P���� d	�����qޕ��A��跗��
Q�88*�l�@PImW��W��-<�z�Ͷ?�E���-a��2�IDG�yTRAOT����h�8�|u)�	��������o�-��!xVo�W7�;ٍ��/���v(���:�p<W���n�$>Y2}�spi������$�6�C\&�<g��C�L1>t��҃v�-�5�C7乲�*T���WD��o�#�l�='��S u�f��b\�a�\�u��5t���_J {���A����j��9�|c�!7��q><��D�:f�Nf�^ �[���j$�t <3��w��9��^�����Ԇ����_'XԖHTv�+�莏��U�[MK�_�YR�N�4�uJy���1��q-7$٫�� y�!c�Rd���Q#��X���GP�����p�
ƞ��0nc]8�j��w&P����ʳ�O�R��V���ۀ��!�z��!+f�?P@����r�[��Dn�X�F���i��0���7EG�R�D3�C8��'a�`��~:+8KHguH���,�,xc!�19&�zS�Mlێk$���\��z�-�sd�?QKS}Pt�>p��	���M���t#v�&�k|Rn_���*~*,(��#��
�k�4�^���)������V�{�`#���-�p�z�����1� v�t1qؓ�I��>m��{CsB^��7Z���]���
�C��J9��t�4�_�}��հ�ة1׫"����N�.���B�Bw�#�J��k�Ο�n��x�,�÷�N�E�n摞�P"1Ύd�v�܋�uKߓUv��8&ZO��[?L@�y9�����M��tJ�>�r��ËsHf��7a�ˡB�
��jQC�Y�Ca�� V_��`��5�xM��	�������ƹF�;���y�v����1 SG�L*�L3�w]V"��w�3Ǫ��I�\*fJs���9L�?ͧr�{�G�X���	)�R�XHrreiC�j���M;|�C��.�C�0
�Ҝ���"�\Ѻ˺�qL�i��r�2dMX���X�X�� �x���q�YN�T�{#)��O��@\	`+"I�r2�6&P^ѝ��_i�H�v�M���K�#r��Ivq�#!�^!��	2l��
Je"��0٧�����X��"���4�&��\b7�����z*P'i4<'X0�8u�'�:��HlA窊D���v�!�P>
���k��b[Q�������;�C�q�+/�mC����T#��*R�CprSE���1�ݙo俥��B�̘��*2��9G���2}�ϭ����{;�u��%9| W�U-!/����A4�qظT=l3
�ם�AV1�p޵�Q�`���� ��9pǱ�ͱc ��9x#�H��h�}j�Z�U�i%�$�9%�9��D���f��J'�3��Y���>�)���L�!��9���M�z�.�lZx~B���t��m�ꉘ�>���H� �l��0=wi��S�/��]�#����2��4~z����ʟ �x&
�Zw�U�&�ޜ��L�֌��ͷ�~������Y����V�l���I+������4&������.:��nn��3\ۨ(?�S<��ۏ�tv�s��+�h��k��DMt�K͟����>�-`�|�zH'ccߧ+72����1F�Q�I��()��X��5l�g��mh\%:U�
��W~1���o��~��j�|