��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su˸Y��'��d�Ay~�`�i���o3 1&����1\T�����	��!mF��
��\�ݘ�#X4|'�~a	N�1�""rϗ��?���ݝ��^��lt����d�k>O@�0�#/���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+����=n� Lv���:>CQ����̛޺�/�,�]C	�/P7SkT��V���0>�܏�.� Ȩ����O�4���;�<��@}9�M����:m��k#9��{"�r�U��k�|-��s���-���}h]�����)��W�O�b1q�u� P�W�d�I!�J,�4v�u��Ѕr��q� [|3̜K-]�ed�0�x�~ʎ���l��`k[��O�I�j�x��F��>HU�;��W�����ƻ ����Sx(�]U�۪F[�I�����Ǵ���I~�Ďx�
�+���CQ���c^G���FU?��,{��a�"�A�c�T��?l�/捉����[U�(�Gi4P=�\�sX��aA�C�e�+�	�(Mu0tUu�Q�:�_g9Ѝ�_�i���b��zi�O\��ު����a	Փ���P��Q�ۭ���1����$�SQZ����/7a�/�	��(r��wJ�AC>����ơ��ZB�~0�����ю�Tm�p��b�6L���}��Ot<?�=��mwI{�݁�me/?�D�Fܘ�҄����@����JwXE� ������2�nI]��O�k����c҉���P��!��h��^��	�;_�x��g�������s;Y���������d���w#�[�i�E�H�ꈏ�'��N�n����f�
�9�t�w���8}��c�-��HIg�Z���m���8	�Uj` �04���`}���IRY4"(�ͺk!��y�tr	�w/� ��Y+��j8�-H�`8�(��'}�j��ɛ�9�9A+�0LҼ����[��ء0��!���Dui�*x���!�|��t�����	P��	���J�Y���mct�v�Y�(t\�v8+l��ksJH��5��iWeu�L�Աp��r�F;��p_�������������(c�}���&�[�27�X�y�Nd���q�>��4��I��"o#O�l���h���H�����H���}��eǢq��q	��ck `R����4��nҞ��ܚ������oFrİ���'U���,��|#��l��U��,2wލ�(F�!.$����ce� s\i�8�Йz���
���6���UA�^�(7��	�/�Sۺ�R;��ڭ͌ (U��#L1=7``����7�;4Bv�Mak�T��.Po�L�����*�C��bՠ��
C�ҍ��t��'5��I�{���qC�Q@a��ւs��S�����:��B �Zr�8���.AG�������f����5}H�!��@>�� �F��h�M�q`��<}��%��}�{���9��D_�Եݘ�xf�y�0�B��X�5.�8��q
:4�6�j��׊#�����z���̈́~�րaG$=&m������g*5G3�*O�kr%�ʶJ��ٖ�~�L���Z
���l�q��s���̬�F�Gasi��
Ý���.G�������Ӆ���F6��"���'��a���VV���(�.s��(�<;F�w,:󢆙��P��Sw@ͮEn�H_��`����It'�Ƴf���@x�V<�_����F%���V{�7�6ai�$U_�����ߞ�62p��`J�&����'�q�7'�x3�<	�"��.:��/�����#�����v_����}̏�0$(�_?�8�o4g{X��EU0�[j�unKE�4ȢS�����[��I�q��T"�K����l���xy��u�H�y�����lXu	Nn����s�����W�;i!X�)�Lj�X��<��[*�N���a���OV\h�sm���g�%�@(o���H9��Wa�c�l������{�_q�s�p�6x����ܹ��4�\>"��_u���TB���De�
Hac p)���M���	�q��X�qc�����D��'�ߞ�D������SahQlTA� ���+w�m����L�i�j�=>�r�ИC5Ss�>�;���k��!�T�`�M֋ј*T�Ͱ/�&�+V�;�惨U�Pe8Y�]!��y��^.��a�e�4��'zq������)T_(^���p-id�4�EjSV���iD�@�.��F�l�ء���!Q&f�%�Fl�ض	���@I%�����>�*h�G�RP6bf|E ���&����\�bc������i@t(��QM:Ui=/���?#B���Sd�u��M��'?!Z6�g����g�maaJ��,���f:�(�opSlW���&Ⴧx�+�3Fh��n�9��j�˷�;�G���L/#;Pc�)~8��5���?�;�*v	�AT��H�;TԊes����oޅ:� ��p/�n �^F� �*B�Y{���?T]��潎�H��^�q|z�2r�L �C��t^����R��tl�����3�S^S�� q��\���ҽ�"F:��ŧ���1,ٲ����Xh��)B������,ޫ�X�Vu ��#��_�t�E��	��a�����#�S]K�-H�\��.ҖP �|è$���V-#*љ6km=�ʦ ��	K�5h�xS.�
�j�t������?�W�c��8�.~\E�:'�d3�Xh)�pz,\�|���B �M�D�u��]]�&U0��h�H.����4g��u:=�]�X�o���f�/�
jC��m�����T���z�B>ɠH ��Le�ɘ�:�$C�"�yK*�9¬JE�:��v�F�{��g����\jA@��}�q�M/�'�Ȝڹ��c]����H�r� ?�zLd��r���h��[@o��-���U�O$v��ցy_尡Ӡm��ozg��]�UuK�sj��Y��74��2�D~�3I��#��`�gc,�4�Ĥ�W�}\�Ί�6��|���'�i�N̍������m�N|F�88eC�_8f��*����b�	�RhTD9�5 �z;�h �ٴ����H�z���;��U.?�����Z�?��e�(��)�Rv�m�(ѩ�w���r�+��6~��f��&3��>1N��x��UNS�����s�QT��	��wXE����ׂ�!��	(�.�-n��Ss�F,z:��n�5��n<��i���Z�]��ݥ�˄�S���)�I�g^B�-���^���Y�j�+�eD%(�fOu�z��w-����']�t!� �cn�m3jO�N���B[&F?�s��j���q������M�i�{o��2
=�� \%De�
$���!�?X�;o�ʤl4�
8r�����:=�����]��{ F�vTq`?�s�m��M���\^w��)��s����A��oj�\Ʀ�X~V��nG���1n���	�	��?-� ���
�N�P���.8q'�rrb�j�L;��e���ve2e祻�$DQδ�N5��t�l'�$�OExG�0�{�-rwO�g�S^��2Ƴ��r�&����:�2���~:��gp�����z�M��NA�b�i�_������A�cD���򔧰�� �hUCNP�R��:�g�L��	�?�C��2��~r���yR�Ǜܻݬ!�&���dx�\����Ա��=���n�Iws�!�N��J�F-�޴V���B���;>���-E�ZC̡`�8��)|�[eJ��ߎ�����8�}O�]�'���U��X.8��	�Ň$�J�a=]9|�q"�M#q�D��\+���Hx��V�Y &BKJ�zl�ў�~�DHO'{1�@�@\iy�zIu�V;�`RNX��\�*gVV$?�e�g_�o��i��yg��4=N����A�Vf��\��cb�D���"�Oa��B&�l~�i�4䎯���+1�B��xR�1��:$�Gt�l?N�+�{S�����;x��m���?~��՝F��u{|pOJ��Nd-��OI7R�ҁ��<��n�z�^u�#��2��
��ؿ՜���I.�N��{)E��f;�!��`�e�Q�Z�y�^����>����f����P���<�Ѭ�u�K�p+�L]fLK���)nNG���C�I��f��|x+���D�������^��&�+q�J!Y�N  e%Z��^����p����͞F ���+���8�w���O{�"�=#����/ǈ�cK��m/��MH�0�B�Nս�^�R�`l�X9� �BΕhN���1�}���G큁P�m�r�dr�C�E>�T(����I!1��t�N���,��֝������v�rNI�P�ҽ�O�摏��K`JoZ�*p$�����6Q�|}Q=���`����_Gv�T��l�a�myN�i����B�L �䔥p�!���A��z�.EN(t��Q��EHI�2�FR-�|W�f�� JL�`\�J��
α�D�q�����r-��TES�B��@Rw�
��KQ ���&�X�1����b���n��ʓ��\��,`�cE5M��6�ܳU� mY���w�|��BO^W�]Ml�S��u�<�b��|�`ޔ�
��d����"a~��E��3��6��'6�L�����bhY Էg	��M5��ha��:�����Y���+U&L���`�҈����.��ё��%�����fb�T]�M�5��q��_+�s�*�t���������0p��!���?��hq;ݰ�ɏ�����Siql�@gY����o��p`r_��HEѦ$�/ݻf�	\'C@p�lx��HF>���k���?���YҴ0@"\��AQ�����]h�Zz�2:�k��Ņ�|� Ju�(����b�ױ��GUeX��姳����-fp_�Gb0Q���H_��-٢\�|�$2�޲߼�в��w�W~��Ů^�J��:�:��SS*M�����]�%��PD� "L�1������B�˗
�D��Ox��:un�����_�Vke��pk����{������$-��L�ՑP��i�N�d �$0Wn����ӫ��� 辎c�.��v*������Һ��.|nBb��,`��Q�.�+K4�r��_�����DRNd�Ч�v>m\��d�ى�@~#�oB�B8��ȁ�}�>:�6�_�d8K���&��q��Aap�sy�EK�S�c�^ڋTM}[�)tVfYv�~Ҩ%��ϯ��~ rwig+x�z+ty+J�g]�i��� �|�
�n�c�տL��	x%������oZenp6�� �f��d�S�t1�=��^<��l4�q��;��{����b���R>���o���}1p#9�E�ΰ+	��a)�5)�;�Y-5{��i1�!�s�z��cE�3�{k�������S� �D�=������Y	g�VX�qO�"�&�x�w+ڦ�j��	�'v���)e��e�r`B	���χ"5mpSY4�pYb�}u4�0��p�T2k���~	S�	b�y?�:����lC�� t���c$���t��/�e1Z���xϹ�&�[���b��Ҡ��l$�7�.���_�oz����"��|(�k;Sj�Y+{O;�ڭ���[�9�Ӄz��^@�
3�����su�]Ըv�;����2��#n|�奋�o}s�Sȿ)��$�P�޺�v�p�!s�OJ'N@��8GϠ(��ѓ�L��E��>P�mtZ+P��ȶ�n<0�7Ibp��y8Br�E4=j�#��Owդ���2D��@�o\Y$>߇<���^dR���}���U�[x|[g�n�mlEL����m�{K�8��XomP�G�1.�O`�	��u�����t@.Er8�cu��wּݴ���v�Kn�4�Ӆ�R?�x�tH_��mZ�(���~�5~w���3�k^or�d��Xi	�&�B�a8V��7���p�����$<�0�%���-(�᱆i֫�H�Y+�㡽yA	,x�9���+iM*��i�Gw�� ���5NxAB��DA3�����6�	��mib;/�[:��E&��{�Q�{���I���GQ� ؀�?�\��NϦ�HE AВ�<�a�H�*X�qk� �2^���禟H2����fTX��*�]��me�Usҕ>��\	P2�[�V�2�\jI��$}l"���d/�q�q���oIM�62���z���R�T��远���Sj|�D���(�jH3���1#`�LHy�O�V��AgKa\�-9�rmv/�{�Z��R�M�3i^)$BS:UiAw��Rwh�$m�Ы 
�N�#t��������]_���F��S@�&ɛ=�L5����Ѷ��Y�լ�QW-Mg,,���X�tX��5-�� G��W$C�9&�5
��X�͚P��є �]7v&O�u@F�Eh��L�7����*.�󏲜���YH$4��Z-��