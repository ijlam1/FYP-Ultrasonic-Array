��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su˸Y��'��d�Ay~�`�i���o3 1&����1\T�����	��!mF��
��\�ݘ�#X4|'�~a	N�1�""rϗ��?���ݝ��^��lt����d�k>O@�0�#/���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�w�tܔ��R�%��«9�;et��:Px�����R��-��CLE nm(T�+�%]>�%@�Ī�9�3L�0>����Q�h�ȸW�LU��R]YB� ����Fù���,մ��c������ �e�~��ؙ�o&�F%%�x��� ݺ���+�RЏ���Rmd��!t�5�3��h�]7�'&- P<=�r"���G]�E����*����fh������}A�c�f��6z�\uV��U��9Y澁�H�30e��,�kww��& �"��B`�\#��B�V�?��-aw���j���*���%�C�Ō��]b�`O4�$�����u{�>*��i�#96�Mָ��sP���P�E�+�wx�+ڸ�`��ɸ��)����ą�<]�+���I7��	�<�:��p���{z�|�x���J�r)�g\C̶7>GK�8i	�
�!���G�*���Cm�!]:Tg��>��zjZ|'uB�?82�3µFt���RJ�0��O�c���jPm/N�v7^+�#O��)g�������l%���֔<R���F��㷺x�4�D1�O
�&*���A�!��X���1� ,<P����[%��B.� �Ɍ���5'�<Dk5�)��o�K6m%��i���v��Х�0�Nt�|T͒�?)�M_ij|O��1FoN�����}��/�4:0QJ�S�7W:�IC������F�����|��l�G�tQ��'E�u��4ZB
���v�7�"�;1v�1�?,���>d�Q#h�(����P�>x��N�ַ�CF�F�
�Y[\9ɖH���C����! �p���"�^l��6��U��,�#�9�=��6,��?�I�9�#�������B	X<Xn�)�XōC8��ﮑVt�A%�+%��a����6er'g�yE�*�,�mu�z��3{������S��\���1�|���= ��qa2&��4��ʀ����7?�lfF�<��GK�B���5�΃��7�E@Gɇ�5�fh_���������$��&آn�&o*v��k�h&�k�(} �R�P��:T#���kO�uQ��70~��@Q�����Y��6	"،,��#�=P]�DA�"PY6Ҍ�W�π�ao"oE�l5`{��bYÝ�k��j��DT���3��g�a���4h2�@:o��=�!�+���g,{!(׀��-_�?�s//R��,&E~�c�{T��dD\:D�lУ�.iy��0ڴ�l�( 1�w3�<o��j���6�g ����\�Q���.�嵈��ַ�gʔ��g�gn7�hWk����,�-�5�,
u�HHpۄk�<��HN���̪��!���$�FI�&������9�O�}[4 ��ls",(���|+͎�7��mH_Am��0A/ꉤ ���5N�MWiA�+�/E��GȢ��c�}�|��z���/))����1�5>f��}�a�,r���R�e[�]��:�ne��Z۝�,<	�7��T�̓@`2�����ͅ���fB��}�´��}��A	�5�!�L%�<Ԡ��3%�'�J��@��utC܂��Z��g�f