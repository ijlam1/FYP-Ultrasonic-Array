��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su˸Y��'��d�Ay~�`�i���o3 1&����1\T�����	��!mF��
��\�ݘ�#X4|'�~a	N�1�""rϗ��?���ݝ��^��lt����d�k>O@�0�#/���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>%��}w�K���e���c��',�s�7u:IҒe�������u�.7������/�����L���!�SH�L�z��4�P��~���Y2xn]R������\_o�Y.���p-A�E�y��]e�R!�zA�@��Q�ט�c�r�Y��Me�����'QN�=�G0P2m��k��Y� �V�ދ��*70�q-m)��A+`���j���5����ou5��%�(>��E�I�̺_�/Nc�\s�w*p��۴]�oR`�%���(Y=�uϫ��5��L��� �aB�⫢�1��8`�\8��t331%�F]�<�`�M,8�zC���+}Q�����eH����DӁᦰw8Y w���3�Aǻ��}�!��p����My�+�@�V�Z��rV��mz��"$��m���Do�i�F�������B���� �O
���r���󱽛,�l� 8Q5�a�䋒0��J�4�:6�.������q�����*iS@�owK�[o�PȀ�Ѐ�����ސ��٦*+(޻%Itv"�U�yB��L�O�^ee)��?O�7�1�m�/�|X�KM�/z���b�*�c_yVƭm��D���H���x��GoAȚ�������c����ۍ:����?92Ӊ��`�.����U�Uv`��2+�X����	Y�Sʎ%�{_]�%h9��WgQ��<Ӏ�z�.���7T�8�]��6ISrNɞ����ӗe�:HE���?�&�G�������\Ybj
��iU�ϧg|��=!�9k��� ���M��MZ�7:���&�<rE�q�(j��ycZ>���	��F�;%-Pm�E�/�b4T��r�z���YS�����v�da��		E7�	 ���M9{�����2�`q[��#6U� Ш�*p*3�	P�'�k�lj���*�%DǢ���b�ӖՌQw24vɋ CP��F�y�E���L���F�XO	?�'+UV�|�]��UJm
���KVҲ�#_��:�<p`	��WZ� �-��6-�qEaO�t�3�����O����|>
�ܸh�Cw�dw�!;.=T��	]��;h� �唥�W��#3�3�ÖoNj�|5dF����9�1(���3�W
6���ތr��p�^d)si�2N�|%z�1DDWe�Ka��t�u� �����̅����L�~LO��K?���?��C�i
�$�^?�r�T�տy7�x����G��O���=KS�
�@��%~�HyR��n�:�u�L�%'Fde̳-rQK����t�@n��7�Cn|�F�Ϸ'o�c�Y(tlt8?z��Ak�b�&����������g��c4*g�;��Ŵ2���$�+=�!�s����c�/C%��7��8<�'�����z����8B�DUʰ����y�U�+��cjB�R����ⲹ�=K�s�7�a�[��0hy;S�Ԃដ#4jV�)',;n���L����h��b�,BA����6��rR�1����3|r��1��%��@���j@�_�n��S�E��$�pv~�p{��R�������@�}��v���yCFXގ��I�/&��(���lI����N������j�#/l����f$
	�B2�ٛ��>��"Fq���;2{ ����0j�����e�5z��=�m~�f�B�H�����k��x��J��.�om�A#���t"!�h��iJL���kif��Q��myC|s�!���)�I��*.���~����W�h�P���F�ұ���jb�+��A�!SY�I9�`CX uW�ڇĊ�����Z�ܠ��n����zf
� � AȢ~�{��;f��?}{��Tj4��[�أ���íQ�)0&:	9���u��?��wrNUy�NЂ�G2�N<F ) =v=9I �6�!<�_f��y$W��5��*���2�.J���TM�a�Y��7~�v�Tc|�i��f9�t��&�`��J2�R��b�'����*Z�����a�!(�ǤPA"n�}�O��u �ꆏ]�9�褢�y䫣�F�GZA�իB^����9�r���a����B���U$iH�#�V�V�mm�B[�"����,��MW��p���*V�� WwZ';��˽�
=CMo#hں��Q�"]o�+��>3�;X�@����
Xq�UV�ڮ]�DB�o����:��h���{�����7q����`�q�O|��3��i=��L�n��7�:ł����D:{�K�7�s7�|E��n�V����*!g���a� ��j��@�\�'ͅM!C"�wo-wc癭Ѳԇ�����aC�Q5���޽�#	F�v�$��;`8{-����VN8)>� g�$��w+>�7�8���ܬ3 �8U���xQ-����_D�}�����R5׼�X��\�������m�oi˙8�Kz�K\�ect�"�Y�a�f�����Ěu����l�U�k�n��,LJ����¯4�=lU�D�e������Y1F�s+m��$P����f8�H`�!:�| ԏO����r�7�=�(�Ұ��B.$���#�5Ƹ�**����#X\ ��
�ҋZ:.���+���ض����w1"����]][ˣ�&_�9�Ye����D���̲�_�"K���������	9�H�����*I#�%9y�}��-���86S������=#vX�_+�"�H��8}�f
��,>��ea�A��P-���Az����ְVrZi��)���ם%���j}\��P��|�������
��hE}��R�,Z������U����ـ��#G����G!�sw���z�rT�L�9��1W��W������c��fw5�dwW�xh
̏��5�!+�T��%��`�H֏�,�]�۲
����b|e@].U�^4n�Y�ef����e��ԔŘ0?}�g��s�B�j �X��2Y���Et�D�d��s��V�`p|�d��X75�F�19�j�g�#�XXU֡W�����B���8O��8�:�̬}r/��zf���f��0��g�$�;�󴚇T"<X�~h�8�(�ur�� �}sYґ�kNg�!^u��i\+�::�'�О������_Ĵæ�W�&r�8�Y�Dؑ�@�j kQ��Ɇg����;^�c=�y�֨��dм�!up���A6�Uh{(aw��`i�/M��#G�����¦�3���Z�Z���6.�噗k���9b,t��S�����8������a>�BH##�~	U���N?�1�6ȡ|��B����bv���p0;�zGB3���y�b]@�eK��!|��� [t�d�A�K�tS��ˮ?P�%��_�"��,%��z��t_�)(z$:���뤷 �>�
�Hh-4P/���7��p*t��rM(��E s��}>��ָ�`�e�Gs���`�������І�
��3�D��b\��A��ʺa�e�)��;�0Fw=�%5�;*�!t*H����Yn\]2��+[T��,�r��B�֩Z��B9��!怈�wX����� �1�c�}3F.GG�}��|Nmf�	+u�oT�nĦͿ�B&Z��_x�!�/�l��v��������N[C�ќF��K�l�w$��jaS�׿KI"G��S�84��<+�¯�<v�Cԏ�)#G?�}�rk*� �q�d�
���Qݢ*����ܷ>$m#���Вq� �Qr�v�V�	����di9I���@�,�����e��wJ×� Ҵ	��@>���N��Ħ�0��y� S�)�/1�(�՝?�b�b�0�H���]ɘ�q�&ʫ�X�'�G�VD��|Z�SW�m��
s��CB�Xy�b����K|�h�����FE��JxW�|�7�aq�H��hJ��w�:��
��Y���Շ���0#̸	��?����������I��RB��!&^��%#9n\j(/F�y>�3��s�߉$-I`:�����=��k��R�������a�4A?������:q$ܙ 1=;[�[R���%[��6�u����[��|n�b�D�8Rb��=�p~M)����>Q��z56�fY�Q�VCȟȩ\oT�7�Ni��0=��cS�'K@t�|��̋��cAv� ���֢Σ*��Ω��;+\J����c�_d��\q�d�
�%�������(�Н�����Ӂ�]3λ.��b�r^�w5/#�P��H��J!"SJOK�j[�%cY8zX�=�	�$"�v�x�息NO��y�;��	vf�i6�'E��8�YQ4z�Tz�G�����p��rG��.�TjU��d-h�E��C7�z{`ޚ@bhr�KYC��^�L]
q4��ѻ[^��6��b�%���o�3�v�c{�}�=�T]�Y�C�i�5�ׇu9��%�''���)�)`(O��ӑ��	h�&����C����0��P&�1��ب�"��`�R[7k�&�ݨ"�MJn`=71����M����vV/��Y�Z0,<-��2TR+p�q��C����P�l�����m ǗGC�r�E ��M�d1��}H���һ�%�j��r��!5��&���-n-�u�4q �#PݠĤA=�0z�(�Rh;0p�u�A?"����v�
��g�-G���P��n��.T�l���ϳ�FMm�ld�1#0����+�Q��QM:�c��{Dk�X�8z��РB������Z��w�E���[��}�M	�,��0�EaTb8.����d����To<�HH��a��>K��Ĭ{�TpB��F�Ί�S�DB���}�[;9�җ������P��5��?�v�����U����'���~vse<�W������x�kX��Q��[1�>��
x�2AKঞ#�B4��@�C�KK�b��C�R���2�k�=y�dn���ŋ5"���^��V���^:P-.ҟ�y'���(�WM�66W�&�҄�1j�H䒈��"���6'�ͷu���E���W�h�"tFP�(�b ���6;;���L��jE��)��_ D���ͦH�)p��[m�=��(_rS:�`(W��*QA�����v��=�#76<�&��`��XUd��J(��pD��Y�6񚴷_� �8 m�Sv{J��S�AU�i�t���指oK�zx5s��X1�-��%&�ݹ��i�U[�$p���$BF-���&sG`�yEM�ϙ9�f�⍅�꘸�'d"����������g��U�s����a�}�$���Eά�-�*w��À�pE'�><:�K�t3���H��d�F�u�sy�e��Ԃ^�����(|�� �w���{����[Oq��W�sbu��X-:r=6���&���L������P�޶���c�z�=��P�/\��C�lܓ��d��z ��:R�CK2�=�S��(��I�f���3�9. E�уK.}"��c��S.U�6��[	e������b�53
y�N�c��G�����|[@�/ �'���=�*�e�C���u��c� ��`�#F��)������KB�b�?B���HG}�AT�s�T��i��+��������;h��?���=x�7���i}�?S��r欀�(J�IX�ʛ���3M�����$8��Ǭ����B���QF�u�!^ffD��r������F�VŠ'���rn����|bV=�0���u���4��{Dn(�GP2E�D��|G��;|��}�pj����?h`��N�lQ�u�GJ��M�p�+�۴��
u�	+\Z��%�xE0���攔Ez���r7޼�`�<-�'�1��>�t��
݊���SBck�΄��~� ��.��!�b���I�F��C�ƻa��ˣD2�ؓ�Ul�`�.2�ƕZ����z]>��?Cn�4�X�C�Oeܡp �W���>5uڌ:9!^�>+�D@+�\QN���n�n���Ko.~�$y�/�mCR�m��L%�bT�H��2�� ��CW�O�����V%����zP��sT�r��b E�ψ�d�0|�+��V(<��S	�[�>��	�g�"�XOξ���TgL�oL�'w8Z��e�<��PX!}�6�0Oc��3J��o?Ӽ�x���Q�H�r��5EǨxx/>a�H��45V"�*�e(��˗g��"⋜_�l�guA�T���4ga����
��0X1n
�:���M�^~9��5K]�X�b�%��k�IN��z�s����Br@�k:����%Y崢�DT�������-��]����u�{�5v���q������G{IJ���n�I��Oפ�����Uz���$ii�V�E�=�Ɣ�z!{�T
C��+�p�K�c9<_�A�P���67�-`�#R����8��.0L�o�*��ߒho�?���6�Y+y�o�ͥ$��Ǫ���	��YPs�JX2q2�`���h�}�r�&%�+~���+��3�1�Q%P��3<�Ӥ/��P�01��M��z��v	 +�b!�QIڠ�I��n6�X��޶�W���j�}4�R\<�qG�3�>|��`��ݗ�b�N�πMv�hO���+���}Z�%k�rf)uԠ!��Wo�7��i��/]�Ǹ�ҫ��UMB�ϟЫϕ
�)B���X.�ݩߖ`��	��� M�U��#9s�8c;9Ȇ?�;��p �P�Oخ;� ��7����H�C�vt%��P�D��e�x�;��A�8�\�X�X�Ŗx���kю��{}\"�~H&RJ���k�Ǖu��!�b��5J���[wH1���z��LN���|MB=�ˌ�� h;Q���d^,Ḏ�8d�Jp}���
�1AN�{,��I`[vޘ��~.G�1���eǇ~��M
��~K���u������»o��a�u��VR�����ZZU�J�k��d�/8�K/�}�@ �ŽN���-(6�
V��N���S[(�z� �H�Z��ù��)�&,���<g��G�8���+��?��������<��do㠮�ྊ]��A ',�j̏������AI16��-4�ΜǝT�t����6kF��6L���<m*�a�n�0#SW�u�׻̔ ���l�)�y�ˁ3�TJ+~�Q��s�`ٜ9�A�^)*�55BN��#�f���ҳkg��F��/N�k7�9�۵M���_�$tZ�M+�gq��=g�{��o��7���D~���یF.��)Z=dlsp����_0���O~�GȂ�����m3��o�i�#w�uT�&݊Q�*N����<R���CJ�a-�: �e�O�dс��J]�J�)��X��!�|=�8P�1^.���:K�!�s磈��s�*"<[ϐ���]�Bě��UHԑE�������5�"0�Z�4�T�!�U�X7�c�IW	������M[��f�.@�r2b�W�,�e�M�.@�����/�E�@����\C�����m�R��_��~tDL�{a��S�P�w�[��e� �sFQ+#$�b�-�!���>^he��~k'8ʿ%�f����o��IbYV����z+���cwVCb�����	��������h|�m �^�t*\(�pyu�޶d�]��3v����m��� �u����;KZ�a�����Pd�%�U%h��l$��v�nP
�rяC����1' e���&է��[pK���6ܗ�h����o� G���t�l�9d�2l��@�D�U�pWx���Z���F�,eW�r��Pv�tmVD�N��Go�^#>�I
��4�1���� ���f�"�"b�,;9*�0�im��)X���g\Q�����	�smk^��#�z�%|�m�z��8��|J����	"�>*#J].*{��op�A\}ۡ��c�V'�����ş6�!Q�0SgTLq�4I�'�[I�S[
TZ�Oe�&��@��!�D&�S��ь��_�Aǋ�Ax\D%�p�*�K틾����΅3�J�/�E_��$��`=�E�[����gfjipa�ᤷH��r���81^; ]C&د�"KN����%������A��8�n�/	CNH��R?R/'@���W�m��Сlc9��{�94�CÀ��~g&=�����������m�)_l��#/2�u�����>�	m�ֳ-�F?ֿG<��!|x���p��+�V�Ԟ��P�jAئ,k���<�译&�f�`lL	��F)qp*�4�Q���V{���O�"��i�Y�N>1�/�N��dha�ӐNý �򳪖蜷�Z�v��A������V<���X|���l!�����ȗ�7H���N�(��+!Hq��~�{���?t��&&X�Y%�v�����ՠ�~];O�A�Q��K���@�{f�=���{(�\337
g�8ޫf��cu�&0�aH*�L�g]��u�\~i�{�����+��+�(F=<3�v���&���j�.?���N8��$!^���G��QTL��4mh�r{�<A��Ϡt���k��<G�ʏ<2H���'z ~z�6�&V�r�MV}��g#���#;F|e%ܻ��s�G �&��3��lV�r8�B!w�w��G�ч�<�2����/P2E8�gS� Ԙ|.n��F��J��q��y�V�@v�=��X.N^JC�:{#ړ�k�u��F+��p�����F�^��{uy���-��[ Ҙ'��بl��	t�G�kiD��ى�lH*�b���%�7q|���{ng����5��ف�6���(f�3��X-QV��w��9JO�"QA鄁�_o^]�LWwoH�0���:0A tU���x�����E7��Y]�bd���O��4khP2�����4:](�����mdxd.+�kW4P�'�B������7�;���x���p��BX���r�(�׸�=l�9̊�y�)��"/���%��[��Q��H\��υ�x�6�|-y��C `�}��=e�KC �g��,�d>v@Z���m��i�A��YτT�PvZ6�4F��?�݁H���&�Vlj�4z3��~E�ۓz�b���և������5�}�@e���G90g�AN֢��]���$\I��������
M�j�>����{Un�s�A����ac�1��B���(q�z��|R���ъ�vO?��eҥ@GD�����eZs�o!�EP�6S��Ƃ9\����Hp�pV �o�� s�����ٔH��3��*v7Z牙�a66��:��M�*GA���).Oɉ����D� �e#�c~��
p�pd#�	�p$��G�~�"�v� ����q;�/9��FN|�/:����r��iE���{.��np�,�<�pu��zb �rP�9��݆R^���û���Ð˰�57p�* ���hh_~����a�n��{ӭ�e��2B�n˖24���NA���ʏ]�!jz�!I%�\Y����9���X�B'�0�S��P�6���X�"L��*���Mt��J�Cl]�(����,��T�a�c�\rk{�7V3cC�{�KT;�kH��qE�5M��RN _xM���U{{<ĶW����n�,������֗H����he�ٜ����2�`B6�UK�J;��imq?��yy��O8��>��_�A	�,�������ޒ�O|��(������������=b�Do4�ѱ��y�lw���r"��G~ �lZ��dόW��Tbr��Q#i2t�����^�C�/n��c���J �y#����/\A<�B'_�M��X�˧	Q#�l��Е���&NP_�'��U|UI���Q��I�޽��w(�@a�.J� ���\�1YB��2��R~�'��T�\���`�H����� �ǟ�o�����~}�c��E���U���6䑞�z-硾8�n>�l*�/cW]�X6������*m��h�N<9?P���Mhe*���&z��q�S܆D��~K'oE7��٨(�^'��K��f=��H%0�@�;	�	��+D�B6�]�D�:�6�A6B������O���9���߸��u���>�4=�--7��Tb"R����A^����\z����N�k@�X��#����:*[��`�㇉L��z@j/�Ҳ�:�-`�X�\-U���q:�2�F����6���ւ��:�щ=�;K�'��Mp��*bǡ��BZ����TG�<��@�>N���Q9���nfŵ[�6*N�mj?�a(���5	�7*��3�ŝ�A������l��f)]PD�'�8�iJ�N�TS����~������D�A��e6���Q�KL\D���(��(����uF�2S����8?��Q���Ҁa�ۆ��"�a�q��~T�U���އ�zШk����-�G?<�)to�(1�d����a��Z�u��pU���S�F�]���K�4��k��VK�&5̆�f�!P��N;�ef�;b� ���9]�
^R)(������M�c.+����Z�z�y(��5C�_��95�%�yx�U��l.�	��X�ը�	�o�U�s2 cq��h�HRӬ��P`9R�$zl�tf/^�>��<�*m�E!L*��E���ۃ�j1�)-�U����F�DN��$s.�e0 ���H������׀�$�����J�F�ܥs%f�����ٺc�52
8~4��{,CV�H��0�g.3�6�<��@��cQ�xPDx|7�d@N5�mW(c�L)N=E1Z��e�!���[��s0"EA5�U4P)�f]�����þ����ٶAZ:8s�dr��4ٶ�=L&잻偷	� �죈��v��^,/�CI��~�a��K�g�I��x1(�	A�����.2ų�!�����TC��L���$f�F<k����G��P�1
�5�� cr��!�����Tɕ:ZGl��
rB�$ɪ�>��
�I;�9g�5k�� �����a�
wB�P��ry��h6Dn����$Ѳ��`��L*��l�Gr��ݕ��44��K��u�U�@�ޕak޳�َo@����1a��`#�n��g��%Q={Z$i��ދE�b�Ly 6�	s�?r9��Z���.��k�[&hXdX��4v�32��mF�'�gm��^h ���t$�z��&���*J��tZ'����4�O��>���g	e��?N_�IT ,E3�2�Y'�y�`�JV���G"{��d�5�#���}�DjW.@�hPi�ݗ_UHh�10'���=��Lh%�@���
����<�������E���kFa>r����
��C���G������ɲ��MiK����Q�@���8����7��ZI�#�&�A	_�o��k�Mg�p�Kʢ��tS�Kw�ي���ZT�c��������}v%S����8/LGڭ���b3�"�7�+]�LLi����d6G�+kze��i���)e{胷Ft���+��