��/  9s%����;��2+��Nk�y$U�c#I����8F)�}0n��q���̷��#q_���|{su˸Y��'��d�Ay~�`�i���o3 1&����1\T�����	��!mF��
��\�ݘ�#X4|'�~a	N�1�""rϗ��?���ݝ��^��lt����d�k>O@�0�#/���J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv '�\��$0kk`�����s���,��K��mn书�6g^$�' $�h^�ZC��Ba��	ҫ۬mL�29U�Tt�u~6��*g������H+ ��?P��w�����k��aL�4_n�[��$^R���S�}c�2������{��q&|��X��V���[���H�ſUuo�Ig�V�x2�e�f�v
�O��<��}J,�8�ǘ�EgV2}�I�U�d�J��,!l,��)�S�8)�P���Nj� Ï��d��s�����&_�ch��Bt枟������hͺ�)m��x�>���D$.��:�Xg�\���R#�@�Ro���SB��u��Ǽ��*p��ôrYj���p2��0���-�E4e���3\ǌ���T�
�ǺM�/�H�Id-�ݭ��*ߤ��3�f��'�+\�P%s��.=�,ve;7�
#��߿�/��d�zt[��9��i�[����'����r��,��-�FsFc D�@�_D�a���F�ؕO��5 �sg����=�W�4<���Dpg6�1C"µ7g舎"P放f$��Uu�_�R[oh�X�i�g��й�,I{r~'}���GfE�a�vAqEuW���<��n3��%�_�a}a89��q�i���v|��Y�VTEI�d�Ά�X�-�k_�S"����Ĺ�Ɉ��%�e����Ю+Y��K��?��/�~<�FH���{4��y�w<	A��`$�;�6$n�U��vnE!�ڗ��1j�a꺍���Ĥ1�)u���C�0�*�+�a���&��;��7���HY#��r<Uy,�ǣ�F�|>=1�\/*E���Ԫt=B�4a��0�c��Ls�~�i_�51�9?�@�h�m���7A
�m"��RqM Q)�s_<����B����]��ej������=�魐��f�-�D�����_AC\ބ�(��%�����@t�E�U��!�M��QNO�Г��*#�tKl�y-s�ƙ�� ��>�ZyO�m���|�}`x(U�۶g�ZF)}�b�Zt���jt��J���*���0�O�D��K}�?�ɠWzO���E}W��r*hf�l���:|9�ѻa�Ǯ
��O�{�MeFU��R����'٤�G�s���䗣Y��?�ÑZj�0M1S&�j~�_ $��ř�d��t�Q�$���a�����z}�����H*�ٗheΦ�6�b��� ��KN,�a���P�>F�K�g.#6��kF��	��C�q[}sL���$���-!��$B�@>�E�v��V[��D��Zu[�!��;Cw1��P� $l�T�p}���5ݱ�)FJ�K�~�� ��%�� �AZ}YD�3q�氳�W�O�i�����=>0����[Ø�RB�#��~�-�hv��v=��J�sJ��]�a �emtTc��B�I��L�vW%,��Kg���Ճ���B��݊)ʈ��0b}23�� =F�E�sӛު�^X��u��B^���;@��0��/@��6`Ǒw���m�_�=��L7�	���/��\��XZ~HQH�7tx���*pV���\��^P�-wV\��K�Z�������F0���mE���{ڲ#��_�gu�x $�H�Ѽ�ULP#�^�Y���3�3T`!��v3&4�B�'f� ��0����r�]sW��`,��Q��`�h�M�>o0f��p&� ��{��M,�Qtu�gVZ�O����m�h�?�n��Nz$P�%��~��	��mPW�"b�Q�W��\���+�.�2��$u����5�J���F�N�z�R��{�"��'J�f�b_�1���
��ԭqԢg0y�#z.���%2���T�m�Qj=q�0��Q�Ư~.r��*�@��x�h��g�>q����),��U�?��!0��ȡ�|M��1��ɬ�����ܷ䀷��S�t�1Vw��P._�d/������������]T�R�s ���"}ۺg����hc�Vr�SrLt@�w�v^�W��B#E���aP���?%��k�<�$�w����8z'H�tfвw�⛅\��Vn���J�a��8���Nub�>���%���@j�fkk�|�[���'��`�B9�ȇ���`�Ϫ,]wc��G���7�����R���Є�L�?)�ąύ��d�u����*���9]���B�d�g��}����D�dY�;�h܆؇L�$)5�8&)��G���w�����4!�2�V<p�<D����m˭�eH�u��/t�'Y�-�!�s�����|��3�7h`�Ȃ�.��
E�L��'	ؐ��g���`�{P�&��q<r0�[��0�,dϯ��i0�W��.K��g&�@�?��h����(�����:V��hbc�!�5#%k� �R��:.�|l���]������r Gc��1+8@H���g�{^��K��L�T;�4o4g/��zo�m�2^M��`�\�������E}p�N��4���P[\^8��dt��񕳝��Q~U#x8��m!�[��[����H�&��
|��G,
�1+$@�m>	ϊ�v�:�d1�d���Ikr�o����y`G%�$4�^m�>�֎ ������	lg~�fK�ARI
��S!³	'G�Ԗs�[(����^�ȣ�8�]���ڡ��% N�k��Ǽ0xD7R�F�{�\��Ԯw���{>�$_1lJ7%�=�L�2�	S�f��S�:w%(r3c�ᆭ@�͉H�˘��V����a�v$0q2s�ƕ)��1�8��1�$�#)�U��N(],[��5>mY�&�#�WbzB����r(��g�����E^�Q���C;Q/نtc��k'A-Ժ5��I8!�/nz.G+ǲ$OSc&C�⁳U��4 ,�m��c���~�g��ㄩ+�X�Ůˉ��-ײHR;P��r}���'4��%{�V�:K ס+x4A(z�1���UH�eʟg�W���y���MC���sB�7q;�ƛξq&��������G5�ml�,������b0�����lXyI 8�id���Ɯ0*�N�Lf ����~���i�@�MUc���B�c�ԑ�l�:��6���nyz�<�|Z#�`�	@}`9ه�v�H�BF��Q��j�3m*Cg�'���́�����4�`ìփ;��݊�s��Dq���:<f�;���E.�r���U�0�|�]�ް�4�0�Za��v����C��w-b����^JbN2y����T���4��)m�)4���9WWA�E>ʴ,q]R@��tv�{���;8���sd�}��V��td�ا�n����O�&�T�ؔe%�(�8�0n������|�Q|'4Z�&<�����S�G���؏���>Ȼz�ۡo���^CX��]�}K��hZε=��#���߬�&	�~ _�e��s$H	�hI\�0���U��1 ~?��O�(m1\��ZuP��,(��~T)���;�.�c7u�w�Y�b�0&O.��ώ�r��X�7.����nȾ��噃�:����w��Iu,�D.t2|�3�hXs���_GR��81��a���M7;�s�{f�����s~�c�ȿP�Y+�l��6���h�S6�x�ݨ5u���9N���a*D�d�&�	�w6��I{�Q���N�8C�)0ğl�
=�O�||ǚ�v]�m�u?~s��eT����������TKsL�W�P��XS��M̩���k� }A��T��Р�z�~�C�B��,����#�l���W�,�*�q�X&�#�Gg^S��Y�yJ-Ȏ��kĉ4�0i�$o$jF��R���=e'Q˦�)vV��K@Q�6r3C���y�5=�lg�y�T�@X>�Q� [tȐ���|j���=��^u��b�Da� /V`
�\���*G��	�Lϓ��C�T�?�6�'̕�$��s��׵�����GC�1��`��p]f��%�*�yd!���U�b+n��?Pc�o����R4��G�y���gt���Q<M��;<����t@�7�b@�Zp|5EdX�:���zʘ��4�!m ��.z���b7���q�
���J�B'�ЂF�ts�w���;��KX}�v�m����{+����!�nUN3�]T��豓��K;�is �h属d��)s�Y�RA~(��ѣ�:���4�"��%�� ����<EZHdiH�(���̆���ɡ�Ҧ�{'�w�.D�'�Y7jP�{׸(A�<��%{���wH�~2�KW~�X���G��l�]m#8&�~�����{u60GQD�ɷ�����@&��o\��J$[�J,�W�o"�g_��Yr`V�J�6'b[H�>P^�"�	x�`�`H���2�+@^�ګ�*���S]!�(�plOVE��"�W��{��rxl�V�e�KP�p^����9q�u��.M��t児��n�0�'��L�T�	�i�~x뒔Ͽ1����^��_�F�-��я"H��a5ִYbֽ�F<hP-$'f���kkN����p��n�
t l-��1���i�@i͝B��ݰ�T(y#~��k9��.l�*!��`$Q��}�}�.��<�����$Gz|���8��l���Yh��zM��#�A���G$�M�T����y@;d����&��竛Ыd}�:�8��A��cJoK���&��Rb�K�"~k�ŶS��`MvbԵ��ݵ����/��{W�E�k1�Y�_�O��Җ)�b��q����XhzƓ�����7��l�oO8&B�8b�����Vb��)4���.+I�q�iA39��G5�N���9ē�{����]�_?:�z�Y����5x�J�sն m�v*�ߣ���X�_h{�8N��11��I�������i���9}��I���u�f�a<\2�8t܌`������C�x�
CMQ���9P0<-�%��������L����Z�ƾ3��T)��>�� =�(h��In���;s�Gѽ �~/UHYՈ_�$	��K#�yF�C4�� �c����
xp���Ύ�F.f���H.DPV�g�n5�Y9*k�5��O&�[&�R�<���mi�0�l�zz�_�*���e�i�fVw;��,�a`?�k�8�9R�[ �?z��]ġ��#���-P��$�Ҫ:�?��Ó��7p����:?_�Rs�Dđ�èԨ�b�����䠾��'ɛذ%���XX�S%\C���,!	S322@�)6��*wBX9�_��$⼸��>�5�Sߨ��:���m�c(kI����׊�R�� a��Q�c�����*�C�1�J
�^�o��>���Q��H�10�b��sO����Sf�`'���	����тh�j����T`�,�a<(r�Y����o�@@I�@$'����ゅv����O2�)�|U:��<`*��R�������ֻ�qF%U@倽������.?B�ڪ����,f#�1��[���;�	��S���`SKo�Ȓ�/fh�*.�Ǚ�B�$	90M<�G�}�5HI�|�ގV<��O��$�Y.b�Y�"V�w��&�����o���5h��������%��`Y�hC�X���B�\��є��2�p����2��J����aX1�I�\6��,��@C.wxE8L��۪g�c����9X�[@�=#�ݻ���@�ы�)k�7����;��rN�B�[J��U� ��t�)������&�h�ꋵ�~[%l*C
���^�佟T��`G܂ls���Ew�����Tf�úr�_ƭީ�Uqݮ�Iz��c�wk�'����JEV�ֳ!��y�9؅�2F���|�:X��&��#���:E�����dFԤ�#�&u��m���vMq8X��	$�˟μη^r�]z�=�"�R�-zo�*�!��Έ�i�
ܯQBj�=�������h�J6i�R�/�<��N����/P�/v$�'-�2��>E��yJ\:��9j����6��Z:�`�J��a@y'��Z=�M/�	��@�yoa^����6����Zg���QD&�|-�đW�3����pk��5}F�6njr���.�l�)��b�!�/8Y�6�.�V�������c'�SO�Zo�1i�P+u�UL�ށ_��W�m.8 (�����	�יݫnzS ���[�V.����	�0�Dp��(�og[�B�]�Y�x��Z��+������n$m�U���2}�q�ǞH����m=����3��G���|�m�GO�(;�a���|�=�8ۘA�m}��N���_�h�Oo�r�H٨�����3���-w�
ᒆ��Ȃ�2�iCŋ�X�3L�[�'��밒����z��`���bzx��:TB[4ě���h�׷��S� ��[vu+_%��`��șq˯��yYg��L�A�A��� �(��i�d+󬣸��X�`4S����?DWwBh�glht�(9�)�}	<ː����'I4�Y7��&ZA�W$b���+�"3;��r���쥍8q���{G%-��'Qy��y
��P�`������ �i���{�O��΍��
4���t���D;8�yTx�
h2�%��,v��V��?5ROM�е��&C{�b�۸�܏�[�Ei��6� |�����n	��OHn���۔�P�o%�+P�2;�)2e؈<��a�~F�a�w��-�{�H �|p��C�iO8�#x'2�x���2N��+��t���K�Eq�QS�w�F�ŏtF�j���CxA�Y'ovk����WEv��ܝ *9cv��="���F���>aAD�X�k�f��0��� 3�$��_߬^���'~&�:|�&�������F�o�Ur��x��}�I> ��X��=��L
<l&ctF�)T�	����T�s�X�--M�a��L��e)Eu=%2˝��Yƙ�A�{�i�����;�lJR���7�<�g����(iվ�u�'�2���ƕ������}m�c#t�?��2Ya�Ԗg�-�	~�h�����u֖�)���m1I�=E&��RP�� )l%H=7��o�M�k��|��W�����N6�Z�n_+�dsa�0_�)C�S�N"^��������W
������]���-�&�L�7�9����+,WCJ��Т~d�8Zf�??��ฉe�7P��͍��t<X�JB1���CtR+�6Ԏ�+w(�S:�A�&H�(I�"��K��x�|_g������1���o��k^�;¼�A*8�[%n�B׎~�EB�d(x"�<���R��\��3+�7 h��
��=J%%�SiS����紻�r�x�D*�F�u��>��ݟT��N�X��s��`�!�xDÝ{���6g\J9O�������3p��!Vg�����t��'��Ǡ�1��a��B_?ٸǶm���i<J�4���!�t�OѫF���@.���!EBg�G���E�ۇ�6��L,��MQ`�*�;���n�p�"+:��O��pju��l����. ��Ђ�C	̐�t���ߐ������WŌ[G'p���`z�%�anPM�=]I���@�M��,>~���{��jϋ���u�ʻJuX9���k	ŷ��R���$wg���t��T��\��*�v���L����e6򶢻�h�:�lZ�i�VN��覨p �3���Uҵ�:T�>n����m��L��d���_���O��@a�qi}<)����fnw��'p��������|:��i���,٨��ѧQ��"��,�;v�~oFѨ��m�n>pjU��FO�z6��i�d�d�Vw�/���[Ϭ4ٿ���K�����OId) �da�ɍ���k"�����`6D̤P8��?��U7�Cx���b���� �)�:(���XL,(�xr0�q력MJ�(�aD5���� �a��cn���}x�+ʓt-�)��8@(�\����xLI۔O���HѬUaLwJC�@���ت��M>�8���R�EA�_+A&��a�	���}˅s�	�Y^_Y@\53{������c��\�ӅQ����e��Zk�p�J���h��_�Q6�����ڟ!�g��3�F)?��<��/�Mn���ܘ3:o�t��k;����{�͍���wIWI�#H!�ӛK+8z rV���t-0��*���XbhMV��*���ɴi��������z��1n���*�S���� �G���F�	�H�}�)�b�tIX�*����>m���:�����:b���߯��zt�|�sߣ�]��M�9��?��9r�9+@���1	ﮈ��\8��Ț�KYVElWt�@����SB�s����FЍ�e��/�_���S@�z(�F��iB�� ���u=A#�Ok���~������l`E�W
K:ғSؖ	7D��[��Ev/�*�d"R��ƛ�o���_7@C"p�����Q(�Yc�D�3�]݇ߢj�������"l��!L�5�M�5��3�F���IZ����<��G��NŕN�k�����ĺ��qξݫ�7�˟�8o�y���@(r����V& ˢl5.{�*�|���C��{����^��3������ml�"��]!�xE(��·�o�٦��Ś�@�Nk��H<��r�#�ȧc�;�[�≖��M͙�e�{ܱ���\2]@@k3���,W>UKv����GW�t���ӳV��E�#�<����wބ�nR�e�S=��Tek�2n�)'�YܠR��v�������-o�qf/hٴ߽�ɼL��+n�a���A3�o5���B�eм}.w4v�ͥ\�ϕĘ����.Tq ����i�`���̓4�O���]QS�7�P�٭󠪞|��6R�\d�&�UQp�F��E�a��6N�@lUX)�Խ���[�I�A��q6
}.i�++aҥ.����:����hZ/γ�QVu_��ZP���Spu���NZ�D��vȺl������߇�(���Q�uu� ��:�M ?Vq�%��_���7f�C���
{�����34����m��^�o���xG��\w���!� Կ`�qv�)/0ow_;���Ɲ��Ru�j>s�3����H@ �l7)�)�D�� ��:�m����Ȁ�H�{�=����L����f�іӈH嬳�T0�cdˇ��/kTat��=� �{��/r��8�(iա����^f��G���+"�6�I|G]I�׏��{�m�#d	q������ $�id����5�3ׯ̯D� �Tc��W/�� �t�0�K��bh���^F,�ۨx2X�DԱw��*��>[�Ac���ܹ,HԔ��X�?�K݌.q�St���ӖA=��:8;H����v�
��M��;�y��5x��Z
A�.T�e�Җ��#�AB�o�q���!����}	v-體�2*J׬h��ij$g�:n�M^J~�X�d|�.�
�Aw����?8��)}��#�)fސXVx1q,�ĩ:��zWԎ��x�qP�uŊ;�'��MN�q�r��=%�g3�3�X9� �|��cAw���k����"��V���y��,�M�ԯس�$���M`�¶�+�(�j}O�
FR���L�J6ǡ �"l�J_���v;B�J+������w1��"tI����v<�F�`��^wlX��4�aĴ��]�$<��	 �"�Y��ڊK�7�7��YӰ	a�~�9K�ޓ�Lk��e��xwJ�*1��b��v{2O[m?�n1G� 7VZV�"��d(?�������ҿN��%��1�Iq�{�:"��)��'�fox�z.�@�Z@-�Uݫ�w݉b�n�7�g�b�<�:�q*6�pXF	4���-:��u��J��f�]Gћ�4Z�Sw�����sJFS�d"���ofKL�<w��Ou%�X�j�6GW�=3����hp��8�u��ɹ�6=��zD.�ߣ�o�Gg��Jm*̙`X���0"{r���������*��*�݆=U6�YΖA�>P�0�{��v5�j���T�F���}djw�C�:b�.{.ɐ& ��}�+'!J�p���m�UVrn:��MxA_�R&��x���z�'�c^�h	4�/��}��OI��(�xg"�F���]�J� Wt|�z�h�?I˥��#�k�j�z(��Ǟ��Ɋ��@�y��Ė��͎r#i~JS��x�>(�ʸ����������a���ձbh�~0��#H�3��&�CK�7]�I��8�Az�&�_"�L�f� ׍`A >;E(�?��w��E�S�L"�N�13��؀��5<:�����)���#��#�GG�P�&x�=�d�1<�9N�إ&lՁ-�
\-�i�~��%��/};/�b�����ƞ�,��B��������X 	[��&�ِ�ml��x3c��R����vsݲ�x�۸� �"4�$��g��&@�K��	FO;�J�P���ۊQ�m	��_ B��d~��q��\��@Q�E���.'�9Έ[tgx$(��A�n݋��ޫ�N�\,k��>'s@p[�v;Ш�,#��,���:�ߤq����Z3R����Rc�vX\_ ��_�#��"2�������n.xn��7�������꺄���|$�r�r�G�K���q��L:�����(�� ��.n�@�U`4�\j3�n��W&�+���`~
�i���k��փ2_M��O0￫d=S�f�>���5�0�[����ڬi��*�ڣ��]4>$��������KՆh��>u�
�BR���<����Ѱ�%;��~�g�y�M�<{��R�c�b�+�3��PEt�&_'s	k-���MX���8}��%u��G�wk2������t+_P��ʥɎ�Yh'�%��2tV�U�I?:!��*}�ӫ���`�n���wI�Y�O+u_��jfU�s�(�RѕH�Ě"2R&&�V3��pq�!	0�P����?�ʖ��a^W�I\m��_�} ���˩r�\&�R�Lm�1}� �h��k���ޖ�a� �����h������?\����XvK|v�����@����!򑨁4��n� �u��D�}��3�qĪtʘC�+jn��߁G+ˑ�v�rt���$H0�JِΩZ������ͦ/sw�L{����7�2�`�9��t��	�ѝ�)3��9�:b�P' �c.$��2}���J`�OE��h��=��<%Y{�9�ǟ��:�4�:sG0pz�>�������9hD+��c :�F$�[P6Ýe<Q��9��?It�2�3�}��`���9~�\U�w��4��b�X̲f)��I�n��D��>�x��L�wE���Ai#�jb#�OH1V����$v��!S�WHϭ����牣C��kv��?�=�S�o�S��q��TT�%a�p=�r�g�G
c���OS}��[���\�o�4�;��@�<���n��
EB'X�qf �dRZ�׌��2�C��}��c�P��K��":ƭ�B
%k���*�'͆��:�W� =��m�$�y�ʺ��~���
I��È�BMU�OM�}j��8�o�������F�Y��{��mB��<��I0�BG����-w���VH��rܝB����������3�h�6S&t?㪶d<� ��b�${Z�K��;/�X�X�ͻ�C��4�O��F��HP�w��e����G�I38h��_�&�:��w4����k�o�P�V�9�<�.���M��ʘ�I�Z�G��O��=jB���G}B�A%&�;I(����eg���d��O�Wf��Z���},���nUd��T��Ɯ'EA��$tϻRX`!s���}x�-�X��t;���t5�yh�C� ��i�i��:J'�*t!�쾢Ҕ��p
��ٵ�e�4�� !��H��g��y�a.�wU1#l��/�%�>��(�{-���`=��^D��A�_�W�h�����_�^okU5�Ѷ5���Ϙ ��.8,��u5�򑖑cc!уߍO�U��2ʃLwAOau�iq� ���I���ByP��/˧��Y�/��~�*bQ(��#�Q�Agꄳ��F��9r�P�=y�P%�l�E$��/���q�1�ʒ��cV5[u����_խ&�!n4���T�Q-"��~��B_���� [�dz�`/��k�w�E.-��d+�Z�$��ߔ���p �R�*�BW�>4(��f[�xR�<�(Ӭ.�l���h�ѿ�Z=,��B��D8�*=PM�3�F'�7Q�M��Kҕ���h��e9�ϯ���9>lͮ[�d�_1Soo�%2�t6��j�J�k�Y��s��fX�x��(,�Rj��#����kz�Q�}My�)#��5�!���د�������U���g=��fn���ى�I�^O��@�Eq��=N	hԢ�+�fp�������1��r`����"��[���M
wdXk�H�j�3��ѼL���Z����=����X�w���q�k�K��M:���!�Q_��`cB�ì���UǚD@L��U�}��l���jV\`4D-)E�?L\�����A\gr�H�q��ڞ�h��.�]v� K�y7��qO��1�aP���,8t�~�Tݼ��1/���#��"mykĖ�fNê��󬇊�	?���Ln�³��x�v��:���g8�:�Uw26�D�y�	%˿Α�J�v���5���贆�<ݼ:m:W��e�72N���4,D����Z`��?v�L��M4TU�\�kQOEh☈L�.�����]
�ǆ���P�:����{TDG3ƻ\�`1x6��Ob�W��n�qț`�t��ͧ�����5姤�(D�gb�E͙�"9 �P�Q���:ǋ�2����٣dx-��g���H��c�Κ-����3�Z|0$��s���D�jZ�d�H��i�k�!$_��zEd�%�1_���U
KA�;�yI�K�{ݒ�"_ٛ�?��*��,;��L�,��ʗ�5�ƻ��(&i��љ5UA��h�����_C�Ә��)�]���!�u���� 0��.��h���n�J��A�9z�Sy�z����x�g�H�J���^�.�����o��Gf�)��H�2Ū��m��.�.���-Ie6d�1���.Q��89����k��V�$�h�i�]��d9'���v�Qu� �T�µ�d�Vɟp	�5d"[�k�����}/�'�Ɣm�*������HY�j�xl�}�bc�ފ��j{���!|���.x@�ֺ�k{ҫ>G�C�bK��%��͗c��)��m��Y�6תd.d���lb]N^���&���8�+W������`6&�Yp��6Ek��q�'>.xe���'���ʗ������6�|g�PT�"��oIv�y�=�����-�&B�A's�F�7�뒘�h]��5��k%l�H�h]��� ��H�ӑ'h��`�[�	�#�@�����p���5�]�_#�"OA�,���M�2���ԍ��DiŔ�6��.�hC�m���/w���x��z1�i?f�X>j]�ʱ�8�̊�+_��rlq	�*�B�r�&�������"���>'�W���Gk~�4�cS7{��PN���V���&|�@�~Dn͆;ڒNK�P�_��}P�)ޱjTY�5��Ȁ�\sj>n+��Ĥ���ߔ,�gfV�[�����_uX�]x}Ϩ�Q
��x5x��(�%p�Q��ջ��)11�|�gT�&��Qm���Uy���Ϭ֊�:Z��j��fw�Y�([{�f�	�E
��1/j�7�X��a�AԳ��N�ϲI�ȗ��t�I4�����q�;����r�JO�G-�̛��5B�2�USoc˾R��|k��>�2]�=d�k�)��ͦ����"�����u���U����q+=�i�Y��V4c&���L�!���'����6揖���X�1ٓ3�����td0�5��(�B�?���Rv���-��L�P�D�Dfk̆�/���]�՗LMc�~n	�ӭ���F#7��qn�,f"�r�~A�5��=��QY�Ϩ|
�K�SK�}dԊ�$N�ݒ;��ң�x���y�ǣJ�Yb��,�D�!׍}%]�dF̂�j-�D�0�H[����?�+�����>ۺ�l.��� n��*���Ef��þŻ�����l��~��>Ɛ�ٮ� �繘S�����즤���ȍz��@��4��x�N�n�fu�m�rV���?l�f�`ܸĚ�3[��3;9V�`������Zڵgғ��6렻�'	��׺)�o��> &�*�#YkP_$���F H�Q���)���/D��J;H��_���U1]���H�e��ѭ�-�#������d<�\���MW���E*����2��=.�`����8��TɌ��Wfa-�[���ǉ�:�t�$���udT��=�9]0�a/z�*�#88'g4�_�M��P�+֝5�t/�'$!�X]�_]؈bFv y�2�����qy�[@���J@����_r݆0l�{�.��V��t�R��}!�poE �x��z�C*$ �aB�Q �t'9���#�(���I�-p�e��ؤ�g��=�e�'lP0y,��ҁ�=|'�_p��1�Mإ�vwר�{V,]��t|�/5�+��|�l�7��?	�P=�%Y�&�� �����y�K�Z����;c�����~EU;��~�տ҈������᫉l�Z�"c�2�M����%�7�3r�,"��N�B!f����L�x~��`"V{�Ր֨�ѽiv�@��W��֦(��Gz���#��i� ڴh����k>�J��9Z�k�����	����_
{��H���v��뮓���u�l��v�F�DK�,�t	#p���)���Hj^�^`��X��`����m�NÐ�2����m��0�t�7���ߐ��)wb�a�Ӛ[sS���F����"GǙ`"�3���)j��'G�߭xڟ�٢r�e-�[j=�6i/ۂ�t�����ɿ��-]&Mzh��(�pyc�S3���Ud3{2"%�&G�)!]����d����6��	w&�s�=�c^fH����/ .*�Vǣ��i�\���d����Nc�'6���.gϣ�k�9��� n-�f"?� ��!�#|V#�{�!H�P��u�>��o1�^+�!����u,ػ�c^�_�IK�#�gT���G:T���b������~��f�KS�G�h�F3Ȋ��O`�`�7uv����@=,,t<���o{��N͞;2�Jaղ�V(2�F�=.�چ��	�k��1˜�k\|����7�?��Ó�oO>ݥ'�q���
g���'�O��=�^UP��{�\~*�3yj��c���b����3� ���ٔ*�7t����WB����b�R �q�,P�������;ϐ���y@W@o)��v�UEԣ<V,��9��Y6%Qp[�X�Q���M�2Iɢ���	Cv�p��J0� {�q��jv�-sye�[�9�#�8�b~yH����_Z�Ŏ����㯠�]�L$���|��� ��ukh��$���5��;Mcq�/�X���2�qa�i�vt�
F�@ ;<�6�>hȦ2�*����i�SsC_�U�Y;��g�]P�}��+ƶ���K'�8M�}�F?��?�AUa��HU�A��eU�su�E���龟6]ܳ�� T��D�L`FbC�I����֐�s��tNPʙ� Z�2��%$��Ze2�0#K��ƥ;�tH�w�p��s�Y��~}Q��D4���Z����:E�*��[�Y0�d�Zu���kk�%�MY��3PdE`y�NL�ż�K��T����Fy�w�����)�}��)��:?���������G[�h���Ͷ�H��(̆�]�+	|� "��ljA��X<���zC8)�n�����q���|��� �q�s��D�l�����^
����>#��m��n�+�eW�| NF�"�u�K��j�,�5��	H���s�a�(�M'E��1(�+�c25h�� $��-:�����'{ϋ���9HБv��8� ����4r��O�L�W�X�'^ B\x�"�<��4\ΦK^�#ضZ�@�$d5>�t�B��\s�Ѧ�<�U�Cu�0���5��"D�Vr���<����xF1ftf�v�Q��nL�-rT��̊[�N�7��=)��c$Pj
��!�0yv�N�K�g��[?��du!M�I��z���J��{xű����/�=u���ɹ�".���,,���"���I7š��aE�j=J�K]�$>�qb�2��N�ͳ7`�TE}nn�v��-��0��PdִpƢX6D�3'b@I`PA��l��E�"�
)���b>�Y���E�M��2#�8̅�X�M�_�[��%x������Wp"���}�Ǫ�j<�*1��rc-:����V;C��"Ip��{�c]��<����`&��cD�R�K�,^���~�iHֳg�:)�Q!-���6�Yk��z�[-W��by<M�@.^=�ܨ)Y��崬���ੑL1=��0J"!�f����)���z�Vw�N�_��R�pv8\�`���L�V@Ɏ����C*|�t0�F{7�&�I~�.2M�� �Q/�*&Q
�[(�i�ҳ�1��h�Q�o��y\U�S".0vHB필tɴ�^�uo�\��
Vo
�&���UY�?Ӎ��ש��+27��th��$�$j{�ۅ�*�8��K�w��f39�t3�
�^�y:�Ù��p�ƃ��]��+/Kܘm�^�S}��n� 1Z��e�6HQ�=(��=Qu�g�Ŏ�����3Wq�vR�X�^�ZxjC�L�ԭ��В�3�،���ؠ��u�p�2�Z'�`���s��I�"�ʮ�г*$e��#�u>X��,���PSsG�Q
��}�c�`��Z�y ?�CM�=� ��*b�5W7�T]רe�-����Jq�v�O;��eb�>X�A�.P+�g�x6Ya��ȿ�4���P� +�b��>Um�b!��,�m"ߋ��7�6M�>R	,�pΐB���tG�6(�xL�ٴ%�����:�~*90��+Z���Y 74�����󸌼9�g��yT+���w_���zK_��u�+�%�'s0��`�"���D/mӧ� ؋Uʝ5�oVV��A�<e�.AC�*;u�?@�%�����w�\uV?�h���"�n�`�L�g��i ���^�	Ŷ��7ھL\�fSJ����8��=ץ�'�n����h>D�Ѿ��E�P��}�[x��0+=˴u��J��f��>��4�rt�h���Ymoɸ)��V�1���O����yk�O'�9M?K�����&T������Ks:oY��I$�Im�=��j�H_��k��B+� �����T�t؆� �ːKl�0�[�r{ƌ�GWH�ݱ�jٗ���C�<Z�n��
;���5���J+��܉=�\�D��݀M�h�a�E"�}&�X?�U�݊Ú�V�C ���X�7�H��K�F�5W��K����F(-ė\��9�=������}&ɨ��>9���˷Z� ��/�oue�R��d����ۓ�:�+�� ��x�G�B����8���)=]M9��ہ���rјm���p�bQ"�o?ݬ[�
�O���������>i&��_ZqZ�-xa�@Ղ��-������C~K)��j��ֽf|�!{5�ɿ��^k�@�Ī$!u���^؆��<�v�w�?�Q���n�Jr�gV�G9�e~�/21�4���ܕU���.����&�ލ4�����.�6\��W�����U��f��#r�W����űqA�+i�v/���v81�L�x0l�ل�����U���9\5�ﳦ��oYS�91f�hc��=���\p�~�ǚF'-��[fͦ�mFx��U��R���r5#$ܕ�������ǉ������+���O�h�(�Idx�8��Ez�C�kE�+]w�e+]S)�i�.5��9��9�킞���]���!���A5�χ�l���L�ӛ�t�g�-��@�ޟ̾�e)���W�+lgQ�a�š��
���~�k��U;�:�����5Es��I�Z,��S�a������C�>@�*�������t��O�p�������"_֭eEJ>'���q���0rVٰ5�F�;�_ΰƱ?��4��9o��ґ,*B� �0'ӉNx�r�۰L���J��CEr�"f֢A,����(�� ��#�y�G�Ѱ�(�9GZ�yӐ_|���gVP�r��O���W.ռ�Uu/;�����'V���g�����oa�cmU�nS���u፛��a-/�b�#���Z�O�Q@.T��O2��� t$�p�5F*��o�ڴyj���wB�g�- �f"���m�/iA�4.��N�]��ib��5+X3�;-x_�b����р?j�X�3�͂����=,U}��xc��́ /sv�&���"�XF�OL�O렸V5*���b'5�=��B�ˎ��ϛNj*�a!>yQ�:X���S����:Q�T��^��:���C�آ��M��	�9~~7�:+E��S�MU¯�^�]r�����>	$�r�E
�tw�r �v����_��ztI�R��=0���+��4�:h*����VJ�ϗ�˦Ji]!2n�����E�	KX3�ӮC�`o�d�Q���p��P�J)P'nC&����]��C����)/��w�m��fФ��T_}��"e�Yag�A�Y�ƹ��f��o���~j��M����cgm=fo�z�n�>�".LBD����-b��Ω/
c�Gxu�V�>����ڋ��O)hM�����MjsV8�@,44��@�g�\��c�J����u�rp�n�`����Ŀ|���HW=���h��1���2+��ZV��Y4��\"u�2?Y�kM��ф|��V�ٰxHʐUǊ\U��q�3�I�
24͌�Jy#�w��	bt�J���Q�`]-�gmD>엻�z��B'�X�zt��R��+c����{��{E-��j�y���@&��h&���cI�i
�r���B�1|u�b�?�g��9Ƒ=6	�5և�uN1Pu�;˭��ח	(�W�J�iF��nO�ViX��|����
G*J^���v�X��_����a�H�%j�[i+Jw�E�1�K_ExK&;��m㘰���	x�D��<H��$nMD�g����h���Sض��l��\6�8����q�!�Y�"��N}�X�@��{��p @̜{<&��T?KY�D1��lnaΘүe_�k�I�}��&�ݡs<�d�QG���	�����ȟ����,�ƙi�8��V$'����S)A��D�G�]���w�PlQ'��rk�8z4����Ŀ���qF�2�V���$��H�^͵���?���K����0ȇ�֘������?��A��xyqE_SQжLR�k����ok��*��;
.�-ZM+�m-������[�]���H�!��L�k{�G��#,Cy��G���㘭Gt00t[��}�^�p�ye'w�>��XO��k��.����r��/)��
B�����Ik��q��3��̦'5ۭe�������W&\���H�V��lD��0w>|�ӿVk�R�.������Q�j�����w�_�!J�|%�y��`��(���OA�b��V\�{y���.KSS����uXǩ��$0�=n������{������"Zb� �[N��ԣ�C�2:)��Z��<v\kYl<�X��K�L��hB<3%�Jw�V!��Fw%T��`/�	�lmBRΛ����='�[�^� O����"'�����άS�'�bq{�8l�M@��"�Fgv7�fҐt᝘���G1���Rȗ�Bv�l��6�J���\9�Vqy���)$�NDߤ�;g�͝�;"Y�X/��0=�� ���;�J�O�R�OX,��X at���4]�D����lplrW6�vK��E��T�yJ_�DyHP��tT��
��@��!MJΎ�vW����2̿H⸡�X��"����c6�G��_&�\i��0B�,;�#���p���MI���	�r�{`u�L�c.��f$V�S�6����a������qt I�c&LA�|�z��E�`�"�OQ�n� ����Q�1\I����19���y_����_���~@V{�����(�4��q*��?�e����=�@�����\�,�e����in%�_��u��|�1Іu�ע⒦0���oS�%�k9�y����L�����8�&{cK��G�{�/)~ʟ?�pi�����Q�6�a�P�����:%=H�JQ���/�<�����P�C��kԃ�?#_ښ8�����n��-#
y�C��"��3(9�����*4���?�wt>e\P��`bD��B��H�u����ߜBZn�C
� ��Ӵgt�V&Y��>�eT�?�V�WƖU���)&�R��6����%�T��!A��^��?�Õ�^�i���
�z��6�)�%�&t��`ф�e���i:'n~q!:n%����p9��5�"�]���W�KE���y�X�Ԛi&4���e
�^��ɼv���?�	U��7MG�q����&A8;˹����f�2-#K\���U���(�*����i����ԑ�3z��x����z-��c�A"߀;�5����|Kp�%"D�6~
��%���e��$qyF����� k�)��O�R�o:�e��\�[��k����Hr�g���`s�nOL=!t5$�z�L|�}�^�$�	���d�@�$키f8em�E!�0�PDf��k�28�&H�|��ch���.��r�gee獧��p�� �Lx%�o�U��v�"���u�$�2�6���B����0�?�$�
]y�bO&�X�����Fi7
�mz��i`�`=p�Ed����'�z��)�"$����.gH+h�M��+�9a������`�1w�����٠/��c��'͢b�	�?M�����1�H��ߞ��5�r���`ĝ���M������Q�VW"�I�T
׭nĄ�璿-���2���]X��y�Ǜ����)A���Fy)�R���-gNa�	T�O� �3�[����v�A���8ui����4�~?�贤�c��c�>7�R�R��y�늵�5�U2�?�?OR��haj�l^���V'�mg��h�TU6y���N88{�|&��c'y��% dG7)��9�0x;G~�BW�6��`� �#K��g����E�Ɵ�~�?�4L%p@b��aI�PBF���@�&H����`�yf�m?9��S��Z�K��!�.�J���pt\ɷ�\�Zx��8��'�V�
�M�<W����tR6��Ͽl�c�w�*��Jˋ�̝�n�)��b��Up?�3���+e�V��P��_�3�O3o��|��W�Zvn4�@�V/t����~2x.B��m���g޴����r�'����0ZԦv˞�{MM4ΝR�^险y8�J�<$�;L{`d�����ח�b]p�T��^���<u���]]K����Y�$��U�$��z3�U�8�<��n�7��E��7Ռ�ݐ��BX;>N�vh��z��L��	 ��;f����%@y���>�Mx�7�_y��r�c8��2�+�f@3������|e���r�.7��;3��VW0g
/�!�ߙ~إF�^Դ��J��i(�,�5w4Ɣt$��VH'Аt<ҍ�C����
zى��.��'��^~[�&�獆���T�����*i�e�0a!�\;�]"�W��"��y,�*��6k�Ƕ�t��'�q��<Xt��Tg$I�|RGGv(ʓL����C+�9TLA�=#���T�ٜ?O�2vcզy�����і�(��>���Y:�{�Ҕ�[s��
��)了�ȍ��W;*���f�Z�Y�a⿅#䝦p7>m��A���HQW�~�j�7���@� ��©k���V�fV�}(�J�@y���v�'F�#�o�6|�1e��Ie�w��$��뛜 ��Q�I��]K��5锌"�A���{-$o�����&��\/8$I5�D����5�6� 8�}���%��9We��� H�(���^�89F�:�	I�{L���[��_l^wǗ(�P�׈�GyP+Z��c�$�ܹ�'^���8Ӷc�_,7Q5ŹVu�Ӿr�����P�Y�Uf���*�Z�}'�)&	l
ab��e1fE��ȓ����>t�M�]�5�1KH�={HV��;����9�)Mtʘ�x�(6���]���#��T��c��#D�?��?�-ro�'��ڲ��`��������)k��*�o�Cq`��bhfe�
j���z����@X�՞�h����lBg<KbIi3"�
Q�Y���K��Pzr�1����k(GK���$�ⱑ�@�y-X�N�B�#K���x�ǜ�{���I��ύ!^����;ĩ�Q���(:VW���L�`����{�#�:��I|
�gq� ��%�
W�I�`�z��}�2%�ՃzT��.qͤ�19��Y�֋�K{\6�\`1ā�ID�+�-�m����R����<�Fɇ�`�D(�ݑ��P��<�